-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UBCntZsG4eV6xLneiI2+h1YqrdinalrK2X+4F6f6SHTfJah8TjlAfDqjso0oZp3zUtXRGJXcS4sw
UPJijFmaBkQzbZWhvJ+fhO9e+EqPSoVksZSl1EUfSc4mE0rslcljpjCWNtZmpabm8AQHyUHF46dx
CEVh24RGboOznG6d8MGF+IHgJtvJuM4Slh99ZOFBxEm2c4l9gbRiMyFIrB9IVk7o/+Cw3u26WtgY
aw1LWAu33EW8Jjj/x/+1h6LPcp/ijk0+CtjKgO/TbioA1JGjlB3+c1OV+DX2YZjRM9USaAxq9MtA
ma5jCRtDZ/YFXRgoAI1gt48nNtd3TV/G1zOdiQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
mtQxwIcMqrAfzl2nfQ32aBQl60osCiluG+A8WREqV9JqsJz/03c2pVpxyWMNF6oi3Zp1KiYcJqco
pcjLTKQdiYWnuX+y2Ah3uAfZ+OSGe30uTFhqPemO+KtGCXyoUMOnEzsS6b0QYWOyodcJBvgYfnVY
3n6y2pbLIAxvWKawETsM/anFi98pUZZZ6A1j3KGNORkx0eq/lQJfmub6NCUZjvvMxZ57fFLYinKt
VQo+L39mNKPOsoRFpDAa3yNC2QykCNq6hOjz/wugm4li7WO1riAhJrTD+H+NPbSm7KETRgI+Vhjz
Qmi061tpHFZXj+99ZAlayFfPXJlF7tlcy0VF/nAUBLQVBNcQubHi0zMnFRs8+TKh1ox80ZfBa5zB
vsiAKvasivZ5AvJN28aHu9g0BvRGVWk5hGEJETrTp3a0MBYrCl7pcUV1SQrhDPJBxzQaibP/PSB7
Pd6i3WgEKzKXVoqDmRA1LXdoQE+yHLaKYgEZd/MXcSB5WBmrtd/YGSLieR4wd0KesuNGvPsjrLLP
RaV89rxObqYUOOOzhhVZnz1mhSffMZyzAEed2WmBdJ9FxWUxaY9YG65s5cUqfhobShV9vO3Ygj36
TEcyyKQ1lBJMl+q7/k6Ougz0i1/lKp7e5AXsSExdiQoVAPCeHw0Ja6d/OwHK9BDny3RWOKB9GbpD
6VIKdhMs5/KvoMGv3LFtc4pAmTJs1VRJsumN45FRfEiogtbY9qoPIJBVV6VYzjUMYg6pYastxFR4
ArNKXmDlByvITGBIbtLl6eWUPTBVS7dPIIJQUOd256Qu/jE1xJBXtYHI5KN9jdP8xy960lJapwo/
Ytvs1ZrJx3KeIBzD1JzVI43cARSFkRuiBaDs2QyrmvzUbJQp1HEkOdCP7h/R8zAYkzy8Dr+xjsEy
nFmo9l/DD1sOa1opKuyOaEjNNse5v6U+5RXwnaRrZNVs2BOxpL6gQfdXjlubMZknTDApbBO198o5
SoG/RVOeAHjIZyBie7j9Gf4h8utZDgg4gjVB+pZTYHpxYeWckjblezaTYImZHAZgGvwsXkVH2JOc
v83EWpRW6f+cqD1b7sfIxCCRV/RoIUCikpZpOAUNjn/f+pwbhNEtFpNnO7gzYTkoslHug3RxqVVG
PZgBMGPY+AibYGN1Y/ILda24pG0ByOcx6tZ6PzwLuYTP2Hl8y8Iqg6pzvk5+K9TLNynSL7KK8/Br
Ga8Kmr2I8rt2oCHdF+kpa+76QmnvNMoHJOyl+oEbTHuTuhE3C2Hfa/3VaUu738F/dchTHDaEFtoo
DBlCEWHRKATjYNTzE7g7gQ5SJfbjWfdL4EH1/SFCElTzSklxgIoJ21I8af/ZiV2bJ9O9ZXVdFO//
4ZNOk9yy9Cn6XnlelagEJI93h5Va3QAMuJK+2hF3Hkz9YD6mZBXyTHDuobT15oUvya8fVGu0g5uT
LvLw23QNK1Yl8HMJxM0mRUrDR0WolVz8yF+5llqjI5mG4Ci/vkXAMPu3jtqKtoMDhh5BZhYXa1rY
3csGTSGRuerkbZt1/Q7kziw5uTZO24WKA6fLlGjymTg3Ij3xhapYKh9B5/i7r/zNKQn4ExJi/EDd
B5b2zeSRn8jTrAk8dRtuimxKm0H9KMImF6dXr9yikPoHDk9566fzjSaCxZ0b3g4qUQ6X4IPGcsY8
0Y017vYUWEw+S0LFczoh7l9Ky2fEh6TH2hrgh5KrYhzzfpyE5cxrK+6agYRC2ZwA3J2PLCit3Jar
NDqXKvXKC7XjliXBa0ROf+BhR0TGHZ6CCbJg7x+xTf2zD+P4SKmJXkIz6Ew4laUGw1NeiSWswOzZ
DyjfiHPxh/yz9N57foG1SgKF81abjXqDJYgeLML/egBw/OcY6GOlR2bcerb4CzVA/MhOpfltb2MA
d48uyyLJXx21v/PvCUQ66zcGxQ5xT5SoiLQsJvfp8RteSxX20CciEaYR5AfPin+tpQU3m6oe3Y4P
kWNAn+D3uEOHY/S2C2qJza+MH9Deo7YNqzq27dXQ/+P18j5XPULAYt1jnHIND2uRKERpKuAwK7ZX
/RpAriiJCF+xlTt/833mi5WJRKL1MaFnTkWAGd9gr1WZgcHqrxPLfQCpVrD51/Jux/hp5tAwVnTi
ULbJl+FfNK2q8qDKA/CGVIWQW7X4zYSEyV3Wm/RamYgdOSbXNuq1eAWDFSvmQakORz7nJ/K7dkM3
zlJ1r3Z06/lZIpeFUJnxYn402XQYyOZtqUslOrHtg9uIovqzl+WsKjM3vnEgo3yIESLIcNiJao2/
h2ZsCTNA+7my6HYOB3QLsB/TFPWVt4kp/SuR4lJm6vz60oD/w/SAOD8cEUIylPV5N5hsFk6BXlsN
4dlcfNBKP+b339lSYvjBZqk7U2p0EWcQLSklC6KfKgSm8nZQD0K6vl5Wky+NnwbEXqHxZ04wt0ma
bpuAC+l/YAxSjjY/4WdEtW/rLjaRc+2t3OjCF1LLLhp/czfSe7geKfTj2oJI/9FXalgL+SeEv/Im
ZGHw3TeQI7ignFXCetbiCyeqTmQIJB2D3F6pVcwcrjMRwJjN1i+aouTQpQ4bgTwsLgYguigFfDWN
zFu/bzblnDHDG3xmAy0eD97Hl8UXbzu2XjMNuy+ZUXZgBA/3uv3AC9t8ZuKSBFX/QJHjFWQeUEPb
HEJlNHVOc6n/6gJBr4dmOcTJpc360LU/CIrkj4xoC+IggVfj1LwlACfEP+T2m4TGr4yJ6DfknNk2
3CrylXegV0aYRZXwCLIOlEU/YTjPVn4Aft1vCy4g5PFUVjq3QYgK9uv50ejoy1ELEh6L8uaXdUzw
zxMb6u4gn6hSglNKRw15alMzCUsymcjhQ5RjflBuAo5j8D2LwfXb+IDpX3r4/S3x5nlPZaYE/0PW
2mrpUJ49tNTDdnsV6qnE8ckSYwvCUD7ZqyvTcCN49kbZj3knSkEcdcLj2o2rXqzEG2I4NjG/mUbs
ARA7Wm1Wq3LcUkWx/djOWDDthUrKa90CjJNo7rsLJuVPRV545ipqs+llb6kA3M+SDWWZ/jqZI/Uc
ksQtvjBoFSk36Mowj4xbu/gYAN4okhidY6S/lJHkxxf2rYnYACg+/fG1K46Zlh8Ls4oB9QUhbyYm
PxVRvuZh72WFGhF3X427rxwHwRC1rAf2n5UpDCXy6S9uJN8meDmzqMAdAKsBgawZwPFSPrr6UhAc
2Ro2nd/31M98htonN1oMwngUHw/usUCFcUBMRN0lFJ4hRoQXuATSgrCv28THABjsTUAlq0TclLet
IvQ8TD8OE5G+pCXFwcX+DBOT4/SGMHE6pT8XgdxJduK/iNVtkpGNhFAw5hRBMELLT2jYt3t28uCS
EfneYXnrdp7YSdPvkvrHRPQozTh4ju1ffyuhnlafWZN6v6JgCzyAYAb06E4kRsmGHOCD+5Iqx1S0
3LsvCiB6L68fVuka3HoaVJ5OVjL0pdGJKnWs9LAGHzUC47OhVIjPzS55yiuW71RkZI8U94QwsidN
ghHO1OnfBjeB5SyaNsr1Sw9uFo13kCE+CyqUaC3moB07ZOv1CMEBB7uIOtsOIb1JEe3XTe0NTR5Y
2OjVB7flNAXgZXOunZe0wv+CiolMWB4proSZvx3unbmjw2tdeRQYLB/U/sNviZraSmwjS9PVVES0
mPhCDpGzQLAnM9uY4r/s1JqPQoVFljTqB2767aijoEgHgJFtUql3Oqm6IQcxUX9hiFUUnxBn72I3
zMaTN4m/i1hsOehOwE0T39zHrRDJa621pX4B3wz/icerP46S79E3yMFEGa71tGssmDQnsObtW+JR
enEJmvKpJHuFABc0zi7sJU9XLJqLxlpykDdoC8uBoNewES7PHUWbHDQKQfQFmEAUbH05tf86D3uA
7WjOzHfNKUwvNs071QhFh/DIc2tNMtdrwOn41Gu6mCoMDtA8ODm7HXypO0DTFnHKKHrZEPQYq1Mg
GgM7V6XRsxDC4zNEDhd5pRnXixef1E1e2eDF8efZ5w/7EDSzOMOS0wmz7eiJ5sK3Sriir4mjw8H2
nVJWEBqjwl9rggL+eyTWhbLIkViIBW0GQ48rHw2l5IQ029UEFUqabneoQKB1GiQkKVXNpXrP7AlZ
21X7SKlVOzLHtn9Pu8hiU9wfoJMtQNpi6Njx8WqFDzHn52NrwbybdBSIvi4PVduA4gkpvUNcEmOj
ku2STbpg3cO4632AFTwPv8Yun+WH8M7PAK5OzlxZ5anjnnwJf8wgPpi16IWWOfU9eQuzBCc+Xkaf
jsQe8Wyok9373bNSVNIanOG+uxa39b87qqMHp/h3iq1930xSXcgRiofr0Z4UKAHPhNQZSJKLpUjo
G7UKKshykG1jP/O+9y5lqkKARRiI+UFrHVs+eS9FTVhWBV1LWAPww0Q+HVhCSgvBRJAg7fTJ3jjX
008EcIt9tYUPwmLVSDCD+ad12E70qBqUHO2Zd4bGpqfBjNfVmYEjIDD/AcXFwSXww6zAN0hfxx+1
MpbzsBSFLd3O8tBVfBPa8v5A3kPjnFro9ZDu7Iu2pmaaQNyvnf6k7/TqUMrFQccRWstA2YdCCI+r
CY6e8gofVxLC6ULe+XNsgKJONL0vMzWUDw7LO5G6Ii1kzzJLFlPnQlqtCxrTQiHXMB2HfrEaUw72
7YsGsCMeKV5NykCURyosMIYLAVXbIH69Vqkqgj2tZi/CawIDcRL6CIUMMBilJjrRr8QcCiHYT8v3
tlsMisarU1R1tdWYGVrjC6DRMghn04odl6yGBxt4fFD47Jeyx++p5CU6NbAibjvLcXnQCopQ/wGo
QilOiuabjgl4se7v21Jq60w3Fj7S+PoCxMtv3xacArJfUwbAopYYqJp+2+emri2YJCbTgKCxeimE
vcKrhbbYIvu1Z6733wBPjzj0Ow6o13Ic9nvhgnLXWxdNhn6JxkuCPypjDNvhBHpc8hT/O7txOWRz
pFtz2gXo88cCpqkClkmHpVU5LJjqvCq4hwlkXr0z2+Nk/4yUa2Lz9aHQnQgpZWdA23Qmr5wok+7G
qVEtwHV5PorxHNR5Y7qHOP5Z4x2QSWU0zYopeRpvI0cA9c7CnwFj7PDYRF/vXuyAesRQQEW/LQGW
teypYhGrM82xv7XHq3HVWQYcYW+MXNrb0mUYs8vtHVbiFImzNNdxiahlYezXQdDyT7CiHIOLzam8
EhH/YaMQph493AjE5Gf94fWCQf7ktokj4NgH0TAvuxIv7NE+GJFSbZomwNAf7TqebxeIDxjw5KkA
DXabCoAASnRFiy2hXPVE63jxYrydWOdqMuAZjK21R7AQHtHhTHUdG9LLz+NABxG7Vu+lhUDHhCDB
v16z3Ck82Yx1vpkMPVYo2/cgyKdX5Y6xQeKLDDME+ZExJwVWNik1jJY+Sqx9b5LRdkcQkaiSLFGC
nHfZS7LLHQgld4aQATeGaxPq2fyJnQ0IOVb7R8JB1rcKr2gHkazLqRk3HtFMmMlPghSb66p8OmPp
CHChT4XOmH9swcEas1xY8zKGWpLMnPKQmkLxrbgd9IkkGxKorhAL6uy2gzZjaDbDcUsc1fD3SDt6
UACZBaAZU7udsxxsyVXaXRaFwy6A6FoGvLrTNQxYTKY2fiGkbYGW4ZcHpdSX0VK8AL8e6Yjf7WJB
OlDnRMwJ+Mfw7KcyEtGumIlWbu5XLN+XIC4cArG1NpQ8xnZefRgchjjzweNvbRQT6bnv+IKiIFOt
h77eFlpUudHIwIX3O1weyecF2PRAYL99BmdMzakOpdDVXocveFO5m7rUp2vVzvl6+O82pnQHVe2v
kGT5kqPZbVPiOXtHnnP7ItRjsUWEenEn8lMk0VECWthWk9qJe8YMvJL1aUaaTs8ehhUum4cw9x7S
gLseehPQEphrNlM+3xU2soerErRpv9AGZb45HtGw1YESxJLCAsmoy1m9I1ZfqZzzHiG/SbJfcikk
DcHPGsi2jNVZunjkUFURcAK0p8W/xBqjqDsC3Al5QQRpmML7rz3br8QAju/Cvs7l5oqXFKk3g9RA
roWXgeHOe9s9z9HcyMZ5IKTXO+Yq9gfXz+eFEXmP3PRvVYhCjigEabZ9uPgCepBiClcNZI3+mB4V
0GjDdkGjlG8cLKYo07k0dmci5ZOJNqbH3voIEv7R4ljopFfh7O585aHrUHZEhG1m8Onm+2MKDv1w
FP9qTNOVLhMvJdZQpuatgbbWHvkrpsRACAoimWZA84EQk3ANAvh+Au/jYE8Mpt3DrPBKVm6O3Yu1
fPw/1es7WH4inoBQRfErN4NAgKtfmg8sScgoVDGFr3YaGvaK4JOosAsp8VLbAkfAL9hJO55aWCmJ
S0wv8+yp89VveggIGh9tQBOEG81h8brEslHNTEW3sZQLwXy589bk8dEiGuXZLHPq47ISioFmfs0N
THMKix8HkMfu9FQyi6Sj0ch/hVQyrnBN1jdRYZ+qLzGssh7Y1CwnqXqc+6mf6sjAvgrKowrR7ApP
V860H6SqHxjnFbfT+MnKXfeQYoKdweopziEjJ0Z8xDeeQKsaen5f2ZdP5FyaxsdW7J14xA4K7/pX
nDaSVqJE0IbkHRmm9RAVV2iNH0XoFBn8u2Yr5wYbOp/VlYP1sQtBvrP7eBLuQdtTNFd2Z1BmR6ZR
VfLzHu+bVpHNmDA1RlzPcCgQH/fIm3dMViAPyQQxaFJuln7uYgWFYq9jE9ljh2MdqrCvUnwsgwpY
wVhUMK9dSeGOrNLTW8cwb0JjIysYoOaAtiqKUW9EvaZOXxOEGrhVsck9s45BupdkZMGJmU9Dz0BX
MQcPfjKJwkDuRjRqWnX8RCY6RhAKVix2mv8pvRjtm1EBjzgkkgVpKm6tXTH/KPDjesnfZBpb/aIS
9L3KcdDPPFng8VCHGaNChorqsnnJ0a8IHD6UUtgMUznPTV28ekt3AdLyJFHY1+MK+juwQK3omzRI
ikWKAETvRtkpyjw9K6ZB1JM7nDWJLh6nJgmYvKR4DMCNtvbHrj5kWul5Uv+sVNiY4NsQAk1syKJr
mdM4ioyImxVd0bOUXU3dgq9ZNzAjjrKXywWUHVHpCkMFy8OG+KocQjztDqpj9wkluVp18FDTNtMJ
5oGmVF814rvTMGeol0jvILjV09h65dWB3X1ehAGyCdPMl0wMFN9oOYQLOU1+BAhmRGNQBnR1810Z
bX/WURDFGrZcyYoDLXE7ObUoIRcJZ1n/c1Oj9fomiYa5Ownv/kTr8nFLTjcceMpK7RFOp/e/2OPn
LSA2e1SLS792MHLmB7rtQ6wdjDKlpdJqOYfjOh3lB2GLNI0GIhn1VVEsRuJUbPF/GIFhtswAK2yk
MFOtjW0tb82hr0CsvxVY+IuLZ+2ipjAf7mDEyBfPnNQnU8ScPczIo/tGnfJeROb5b1PiAYbXPILI
rmUgGOwqrd1HGyPTZuEXaeZoBhmvgpymqtzvbdDD3f/+sfO9ZnTqdQfPc8Prer429NBaFBPJKz5J
Oahi4mRf59jICu2jx2hN76H5qHvPaUK5om42h5t42o1QFdwDUNWCz5w+y720HDKHjE6HuWfLgnU4
jgqJ4YTi7momc03rPTGLbhCHZM3JzUEdwpiG6ra7CDRNC68RDnMvsORZizfKOuL5ObZD7oEYToLO
rMwECdzSOkKvvCJeljvdIb6SVXLXrGDq13XDXRdmGADZTmod+0H+aC0XmyyuJAClQwwG/GOjepA5
Yp6J+Nm0K3vLa81PEN9SfrVWA2osBu6dQKMDob3hlcBLX5Qa0GTZK+Sc7oxdMraLz6O6FHFlSQdu
DXn1PtWkTfoloOANXhqvVtk8RoOmJXt4joAjLRWWphVReeKdogd3VQaxTbmkwiUIn7vdAQ2hYaVQ
8n9RYWh3jhefO5kmLjMFTYY6aWXKfoKcxW1VpGau/QQ1GEl846XQTgqdS4wuO6Cz4YXozQe9aV9b
/EniLULbXP92tWXthB8IjOArZ1FQi4U8j5y5XrfEBnG4CgR+xY7xbarNgdUxGzCQUnrAQYCjdPAb
xiPRcDwJ9jX51fbYwkBiafE7Deq2kX03S+AfHdOI0QqeBCVzSrUN2sil5wpMeLF8wveVGKcnnCdw
lEC7Kk+0TGHbW0hKE8XJw+AasGPPbWRiij/WpfwxFU1D9ufAzpaecnth6B+U3Oyuyuief8KyJjW9
BZU65lHbb0f025LBUpVmWffTjhSAUFG0ZKICvBqnurWtPitH7P5qs4Uruy/urNWUtrvjtMrVv3JS
/EUIQrP3PTXp05jHYeY2u6E4/lB4LjPckoU+parjTRapZBH08NnpeYnw5BiQv1cQ1ewtvcG42/Pt
yBL2wTJaGFPwGiQ97FXKckurpquD0uKgPONVyG/+UCwT4PJiyhy8vjS0XS32KJGs/yG2Ygd9yXdz
8gE4BnLjJFYXsyFJXQcGZOsdIUNuJ2ES1HwcK/s8iuNmi6YWiPBlTu+lLdcKpPKxh0BJJLnoufs5
Eoqw8l/grFFFyF6KJDhZujW303EVX0ah6WSVys2DJnBp0TXYfZSI5+2sl/cklU9Kzd32DmQn/Vbn
8MO2FJAWPJ5fyC5HSQjx3zpPETSL5zWr5Xpc2WB2HbHUs4sAAAhjl281aTC3UR67S98Q+6v3xB2A
Li62c0Rz/5QMsiCOaBCNBm7A9dq9umD4m8kUxaIiysKCzHx6uguSbUSWn9epxDcmll4OrsR4SnzA
a0e+jFUlcgjqarRbpp9emhI/sEXe0RnfJ4NSU5bhQXhDue5gFBx1UoKHmwrLnIev1U83C/qvAz4n
nknreGGcrlCbu7VrJp34ojX0UKK2wq3EEFHY/kFGoL/+bAhq29w02109wZaZQpn7oJPl55qOdzNQ
JUVtKdksvtcL8BDDtrhL85liFWMMmOhIVOvwedU2YbF/n3qBNBWF3KSrJ+2zTN2RhvBcYTvTV2n6
mhBJeU0MY/N8M68s2mR+F+nCa+sHpVeolRt05Nmrksz3uLcpobzK8rAVeWxhNeHr5vziKIvVvXrO
Azpk1Txpalq/a1mrdRqIafzMN91SvFuD1vt5p8NQM/DVu8mvX3tmAMNmd49f0KonTiqWG9d6C5wE
spUgxhwGyK/Rxdl/sBuuEoBvm/w09iCO3VRzeqaHsVzPWqd4/yRJuSSAbLLMRBVc9WzX6pc+31we
aIbhPBysAs+m8wuB1+/mzdjt8meDKOHS2BlyMhhB+jKiVi6KQeEQEA1N9xpH259Pxc6nNqgmgNuR
E8nxe4lbwkMoUfkpBq0vVDqYusiKQDRmH4XSJIqyFV6nlI3SK6BHudfxbsL8SS26GjAr63ikVKIU
NH+QT1DUbt+jpSkMX91TBXRByuZA8ZolJlmiRKupNQD1yJHLQOoiclx1pd8UPiQ9P7TGFs9SAQjw
+a7ciHTu1h/033CvorpGNfHrlLoz5b+uI0LzaAhiXE9I5y9279ResedJzUfnTr2rP5m/tlaxMT+f
7vJ/GYCfBcbhwlCyRQHPUS8mZ1B+JB4CMuXhIQnjyWI+5ouzCK65+sI+Nh3c4ilagcRISXG4iYzw
YG6Zk9SQJWEngzqi7Ff9t//I6h7p0Xokc3Z1DT4ISK7Vv97K7G9oo3PdjRtElZ0qjCUmwVq3Quft
tOojxRVutL9Ez3qwPcy2YJz8m3zilolqZO8LuqCV9yIQw7Gq+02z1gyJFzyMDK3N1glX7vrDr61D
Znu9zFyDWRUGd7mIs4Np4D9zbBEtNkjvIXPMngSiVMNf6cGJWCfmoPDNzx64ODWcF7QFLVukKjXv
hz48fy6nSwUcvsWp80xwlrWwng7/8aTiJXlG/EGfAMcZr0D8J1IluC6YofZXw0S87eHXxGHyEGD7
SNkQn3DsrB4Wk0uUkS5lN/eSYTveJmjmuq6QXrqtU0WkmNBcQ8jgbSaNXL/9aU+gRG7OYI5dVj96
0cg11wvQ7cfATtofik5eml81qa3+phV/XezmavOm1gf7HXVVmxp3+C12+Zd8h23UCZJXbVAxBteS
fK2wjmIe+uM+v3SzphDP4HMI6004ARDFRpwK3LrAhXqui19B9RDihObP9tdURQQlA3xrwwhjE+92
nEWE2ZNvRL8AQ3RlCtCyxs4YS5pU6JJekpYD6RtuBRCWx8hGAov0NqTsSOX8upQPdqFJbgP5tdUa
PxMXTXEHTuE3d2BPYBAGVkaqw/vmulxCU9MKk94LoBRZgKOqRGzjXJQ19s8NQTKEPnuZ3Ackdt3W
rQj8lJFK8VLIf/U5huH1KmVnvQ4L69SzXD8QGWj0VG59L1AU+J5txXKeDJdBFVioXnKEK/mUNb01
fjxCkdrDV4KNooYJmXX1HsJYrJi4HENtnKVqYoMyU/9cc5VgJs9I3i0Qc6hSseFsw78PXbw/TLc9
WVdeEM7js/le2S1BrGSHxbzeen9GBZp6wLurwALwdyNbpgD4IS/aUQyZXjNgop3fH/7FxIgbgjOL
hEX3OXuSuFKie5S6F8EGNFddvp241Xp7OQ9QawtuDQBIP6xQ6926BJ93TUDxFI2fEGTCmEe801kc
jkFLHDgmUkinYN7RrNj4jzQnG9Cb+ADBS9GXKyoJJrply+8CHjqGT3TXUFZLzO58CLlCq7Ctlt88
MzZPtS+3/qibwit1zRaxrdy1Gw43c8weWdwU5ktCZ0xxHzMsk60wBdbfwSdwKynk+vuIdIYCFvBx
/T4JYbKotEdLJYqwZg7Ktp+IpgMC/TQ+X9OoqX/nzSOXxU3nNtYnw9DIsSkrI3HlBSePvNUl6fCq
6MlAmcwXXJ/HnGmpHDwy565S4CuDf2QwnsAf2qY9dVivLctNxppsqejFCkDciTeazZvnaYoRRwiA
AyRhXf501fV9+P2bhBo4nb7C5x0j608WXMGCtbnzKrpEm0/QRE4d8v6jn0R4I+eCsBWbkWd9teUD
MXVw4sY6nHMO/Bn8x2NWtxynRr183zeuGXtGlP55rS06R9GRS6QLaOsy0+QyEy5zdOG7J8pk/c06
yD8egsA7apn4Dd4jrj6BY0d/AT5Yt5Wl+4ir4M+GB3ZTbH8Uczw3iBI1QxrX9WuJPmtidox9C0yy
OBBI5BUUnMnKhjDJHNUrx2VVSp2Q9mmTL5sNGww453N2Qxx1qTOaKWRPiPi9NfGtUkBTfHGiQf63
WqU3x8kp3QZCZpG8DukXHEo0oCKQkQ6iAGSbk1mTqOXk0b11aPg2Zjg22qrNKU3tgd5PvFLIiB0j
EK6qWv+NZS814VlK/yue7PffZU6KXDHI12Y77wB+KX8iJaZmmJ0tOESOxokA46iyzoFz4BXV0wez
lRunhMlQt3WlId0bzRKPgewelyCo62qmnwwZFfDFayS6xwRtLViFaIkywNWRKM9nfebAn+g5w1je
nOY2/gGTQdjbuEBC+KR47ZlJHVS7WciY71IE13ZLMTL/teeTzpwNEICNwRz05q0C36s7OX6OfPyk
7xJmmcyWP3pYV1ruYGTyZ2HJsDsQeglg+oJzMq1TipqI1/UGHL2jBO0uxMW+4AaP9yFHn6MlFYZx
JFoaWXWRNQlM0BoJ8bLnT2UORR/kKgsn+itzDy691J5MeYhF3RrDolMPJEB8kj6GWMAZmPo5HM2E
2j/DdFyEwp4VPbh3PipYCtRpzj0xfuikZ0IzAA5bg7xX/odENY4raqOc6/6Q8tfmyhbRWdekNgVx
PPv6BeJnbsjB5rZRNQOZyuDte+KNpDz1Xo4n1TKGRmw+K+oLuPRhcMZ5NAwEGyQjcLFAMZzhXItX
ZZxxtjoE1k2qCULfBgGVZCUX6MKqYpS6/YAEAVcNmQB1dyLmYLsf5Dotgj50FDYeQYbuKGkXl2AP
YyOgOVMaovvJ4L+2aTG9C4O8Pff4YzOE7jCgs4H9jMz5SzqFputXYuvUf8tA3/iO/Hq8DVxfH6nb
Va3/gmxJLshB95Xr7CD8NbKz1lD4Plly5ZjuL6q7kZFsGA3eyMceDttKl8b2bYgMU/5iUZSzmzav
X640JKSTcTO6UA/6hhw8j8rY7jdH4+aRBd9XgEmhev0jEtoiUFgh3vh3NTSewAs63CEMdk2hYoG5
x/kY/QoKjZXVDHNiFEjCoyPdi8ux7pzSOg5xqYXisWH0d6f5WwZ7wRNiDc8GEtsuUWpnDursOssh
PsACKqfapenQtzmL1Gvg0LJSgHHIRtJ7BeV3l4eMf+fS4LyLnXG2ABqqm5o2b5Q+KxeZFPbCG93L
V4ivOh7vXCyYGFGa82FWUAWrrErD0wBkG40TJ3455MPgwmCP/tstbXrt4HikgDGy/SC/M753Wda1
qiA7I1aq/FKhn1kXsyynxlmZKduAg2g8rPr4PyzOhJyNXzzX4gpqpOnJkhtZFBAF2RVmtjdWhjtD
cFxXrQhZBaQ1IOMsPXmefHKi1oZ6w9Hqn1S6eIJCex5eyHNs+2F/BK6DLjTci7KAhV9jy0W7Mhrm
Xn61cbTZlW4+//trh9J8kDF2HjFNAqBqD3yjBB17bAnq6bIev3mo1WDWGzZExUrlrFfr3S/Sccvs
ir76+qKu47IwAu1+/8UroOeOpzoyqU2oVms/VAq1n2yIV3rKMCdX2Day77385SsqUezGaymQ+1eM
xpxR8IpZg1C+YVBw53bTVde+115TaqkHqwo9Zy22iv1jlq812kwLsHS0RMV5UaKDnEFtLioNXBTq
I6jKYxm1j2zyz0j4hAGlZur/42Bpe+XgJs7kxyKo6hNbMbISqyzSS8uDgFGH3en2lKjXwFHKPr8Z
g2YjM6qtlhFMF1zskirhkHmFqH814iBV+cLJ5kHpATjZsdVUtFIIvuoHY2AO05gPb8AsDdxum8WT
N24JktFlYHP+W7nCVjG8HBrD5j0QriKAH0ksl4qtyxz3mKSTgxwy98rsHa8Z/46GdYo/Tzx5X5Ht
+J6UlxPh09LXe0LboH952k2gAVuP/LjK+b4K4xGUMaK2di8N6pt+Djei4iEwsecJioXXj7PfWFXq
YpaY6wjl09IMIs3IFGk2iFOUBOSOQCAjSd4Ie9JMs+BXLzgOt6ppnWjw6wK6ehbm2w2IJSfd2Hrk
V6zAKF4piWwcOLpgR+GHcpxIycD6fhMmIZuPV/LosHek2clulxMJ+PxKugJ1ZL+3c6YF5Jnk7OeA
11XrFB1cXMbevqOW4LNMZxWOgtjwnVMI3Zs8CD42wX4G1VM561bP4x+jSxb9/BR337Yl1e89wJ/R
ZTdi3wn2twMEJKUPrrPJfJ6lUm69kCgN1kMcIuFUWioAGWNuXyEefUn6nFlg1UzSPX48b/zS99lE
uiBAQjjkYcjS/WSJnLvB9xMngiEnkTWuwhjJp3uKOzzXbg81HNdOTq49DMsCsLtsb4oKpbEI8fJH
7j38XdMvbSj8No3cuIR2Yl+r5BnZIUxl+yz+HN+lFRXrBn+Gl/AvRI12xnR4KbolOkfKw1qNwu7S
ls+qh1dloMFtllEDEMWVS2LT2MEG+hJCM8zHF7kEE39o8T+Do8b86JhBqlgEc83wab9OKU/H6G0j
AFekLxv3nFGe9ot9rK0nvWx3DHoyjj69Bc64hY3meJG51lJEyUpZa4m+D+oh9rfOBwn49uJQcqxs
qe3CDY550XZHIkI7eQ7UGWVykw5e17t+0DAwJq9nWubzSXOAxtNCgInTSo3tpcOIv2m/EPo8H8D9
bn5tYqg98mRQ5sM+giVA/aSONOhXH34XmQWPwACpeAEYuaDgAO8w/VfHk4F9bNFwnhQ3Oj3LBaJV
34Xl3jFNMmT5s45hVz40wb33z/jy2p6PnexVdHOGUTH3axYNeTfa530Gm58UVW/+qwthGfwRJxMf
FeE3CXGj9vCDujzNfmkUyHM2HXqLZ3rMwnJaKLbfsRTnLFEytgawZn7KMFdiL/h9Wtl9/dGoC+7c
8RvY97mGdxuaNAbHBf/TM8rAyy9JLebR/r7ELvXyqDxXHeNWH4iFQhnufabGLH0Bra03Ky8fx8kM
+ZNMm6hIfjtGxcKq01fjgszEQmYJ/3OyNOoM/MCPotOW231D6mhzYXn+jm/jXE/+4vPDhy3QbSB5
Fx2rhV3Nso8YYEx4Yi41Aqz+gA+wxFAn06a7kTfOjGhfgXPuBVlH5aTFyTHIqvvoueXsHjpld956
ou2bMl8ZFfluw96Op0w+dwiJQ+4kvx/rTrgKUVR3HvXU2YrA/YVii7CL6zwdaQkjXa9zntx5gSYX
XTJfmKS0Z+xqZZ7sk0sfmzZZfJXYInyeNZh4njLpBe78J6uQ52gSzz/v1W9zIYHG8mta4p/Q5Wrv
JYRzWTCmekieyc6IAz0t8kRnmba+1CnQ3ZmNR23e9NlQiM+tSRPYHCWwY+wvJ7Y+HbvJJ86D+tVf
LfE8PBkeoJOIq6cKtbhCZLfBTyUVwodjCwv3RYvgKoiamS5Tiwas+XtXD2kMrNFWkjgDCvND3WaS
KNg272AK2xeXms4e94utIR9dFPrCZY3jTH5LTogo5BxsGhjWi/fRfd1sWx+t0sWUuM7SDu5Dcd5l
XZ/xKh6g3+wpoX9fV0U+/otPiw+FhdZyRYcnzMwSKMsbF180H07V2ehBhs/5xZg25X6IOf2B3rMU
u/F1rGQRbuYln+SnVnm2Ns9J36/xETzt50pIYKfqDCY3gqR3U79JcIdAHYbEq5HhqTyjrVksw20Y
bebMt75Frq6GnBD8EO93VG9yXhtxgWBC+jggfYwynXKKBi2FVb704pJwLZm9Pen4OLN2LyIuU+sN
c3r0ewfrqfeaEebBcqDd7B6DbJTxrltn6wnWsPOEIx4mYOMaGIJOmnkqLqKce4GvAsdoyQnB2lUN
ntL8tUBWyDzAPnAyfzRmbG2NuOwl7ch/7cFtH1UeoxLq6G+l610AhX1j4gzGuvBWk1Dca7yjIFL2
hkZYl+5l4eJU7CiSMtXGSyfW4W/QUT1aRo+A8Pn2KmYbVdqk/KwuB9mbJ98ymdwT2NgJLplhnGr/
bY+gOc+MC0ugy3jA6nX2jUqE4JBsjJ/olcGvOu0cw6ps/Vpshkw0eBanT7CR9Uh9PbvmYoKaHhRz
g+uzsw6N4Um7hO+AcT3t44qI04F5cNaw5Ve5Tl7L22EsW73bU+tL9FIPmoxnNvroFZq91y4FrT3L
Iq9oGmmkmtywuKZrW9fR8Ri6fpEE8YNU1A5sYV34vGnYf2dLye0qXKXhAMJf8miM0pVixzoZvXC6
fl1zpQuQZ8GIp1AFbyQjvJSTrOp1HPhEcm2v8EmCMhpLzOr4+n16xJd3z8EgF4ju8dPWgZnehIMB
f5V36aYtbsE+gVh+FJannNyZiGW+SjEJAfXd3vy4+XNzNn9EzBVPKk7kHEBPPHuppun+Ar4tD5Vt
xNrCYTSqHhRzvxPxzQTpztUt/vnKVp1pCE20XcXRQk7IgCSt9mk+c6XgkYH7QCtSZPSKliBSZN7/
eSNgSnwFX/aDaE2qdcW0FFV0Oeiq724M6HZxiIsW5j+OhhgfeWFglJTa9Ep40J+lvTt5ocGNMx31
dCoG/JNMJ5fRX53ssxSadsz673T2iXQ3AcKAY/A/rNP1yDeiAGss03irDE1dPM5DU/uKjhSZS+n1
nQDwP6CZ2x4UPOvT08Dq8JBwpOmVqbQazagKuH36op5mwkY8XcMcvqHxijx1cqJ9dx6ea2QfTvvX
AppR6kHAQhYlqD7QPxOt6t72iuXHVUxyyj+U1cBTpKCNbZMIkU62iiYz0Z75iO5s9xTfdU45J+v7
lDeRQz+dm1uNxJ4G8akO91PVM/P5q9H0w5ac+dsu5xQF+wtgNhT1QrvgXq56WNsqF36c6n4/tOZv
HgjdqSO8Jnj2ePakHApZ1ulvy2Cofqc2tFSzcxkzAa/gh+X3AoNk1BN9tifRkzFW/SgJ9KDFeuvI
zbMkAVuH5IWgbeQnBLPUY0AstXJn6oadrwDBoGfpCAA=
`protect end_protected
