��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���ۯ>����"H�5� !��3Pj0�t��bV½�Z�B����{���^�C5Pγ�U|G�)�>u���_�@�)n�\i9�Om�	M�J/�����=�(��۰~�k��L�n�2�)�5�D"G����=�7����Q3 ?!����ǥq�{�}�0����g������(�"xX��(*�R�	��^�������D��|19�����OO�`�#`a84��Ĝp�!,��b5���4�L{���Q�D�W�U:���E�n��"���i�<�m%����є,y��[A������2���k��C���ơ���ha�A�l#1.��b�W�y8��B�"%P�r%��~�}5.�`���8�3��>b�����g/��G�MX'�l���|��rR�x�b�=yr�މm*"�x-y��<�T�4��ұ!6�Ȃ�,!+�c�%�
W�$[��_�-B��(eCa_;��2�M�=.X�cGZ�����VC�E��s�\~`g�lP�\��� x������9��P�A�ԪZ�[:��BM|�l;fX�ΧlvX��p#�u(&qVԥ4v����᥉��E�e��� ��Kk��ᗵK{V�i�Ĩ��Y�j(^H����d�)�i%�Џ>{�mh�ũ���$	#l
^���v2��#�<����7 Y4�@A��Z���Y���1����Ĉh��
���7z&��:]��#�̶�6_|cv�Cy
��N��������
esgl:��'�҉j���cH�fyǰĎ��&ed
X���m����(���@a��ȞƛV�0�����`M�r<ޢ$��ȞV�/��rs��[�����x43&��5'�Xz�n(��1*no+�Fq�m�`�A@Z�zAD��	�[4��r�pzGP_�=@.�^��chQ�V(̸t�ƽ��>�CSC�%h�D93L)�SU��Rļ��j�`O�̃�6��l�	2b��C��L ����mh�kGŰZ�~.R/��T���T�f�L���Z�vE��	+�h{5}wӍͻdb�v�������[�E�����s1�"��~�
�W:�5����w2�@Q�����ɻ��&n����-}�����m�63��茱;����O7^��Z܃���R΅�I���c���"X�`�!�� �X������,�}����� $ -˝��Z�����
dM���h�46=�Y��tN� Tj��|v*�s�B_Ï���L��Tu-�?�:o�m G�rJ2�=�h6� �t�{�&���=@�q����z����J6���݇g�ࢬ�,�D
�B�'6�.��"��Tݎ�ا�� k�ӧ��򝔇�V9<.�88�K7M^$_7�#�LKBo@�h�r!-�2�������x����?qdY���͞`|��=Ǡ�9�6��LH��`���Xz�����vp	[��/�9Ng��!�̃�����(���!�j\��OӢ��p ���?��h�I�&3������ͽ���o�ķ�S(��뱟��.��@����y��K��Q�4��"o���6��Ĭ�h~�ꤴ���� �͟'���ZK�+��T �6(���M�V1;��N���^=&�����[��#�~Ljl�c��u�΂m�>��NϷ"�T��JÆW�Z��L?aNYQ�e�@��ib�$���}L � Z|���vRÏ��)�ݿu�/�d�}'���
�m�^�@Z��N�J���bc�-�fV�ŐB��R��G$ �%ޙC&H~��v2Uu(����ԐX<`I,��]�����z�{���<���!*7��'�\�-<�"��n+xL��f�>�Y�j�;�>y>j����_f
��p����hP�i��ބ�� �>b��SAߵ��p6����תK}�~.����W�0\&��2�����kV<~�+��s,{Ie����~z���T��Wp���T��<��D"y�[�V%S��k���d���$B��g�.��I[��Ɓ}�1�M>;D�[���1��ʖ67�ڮM���7���"���q�
C�����6���xJM�T�$`��`J���;��9ҟ�ɮ����r$=�O�2�i�~������ժ�������Ư���ޛ5_�t�0ɍ^< ��&�t3,�{�B �-?%��=����e���rq��H0�!=r�����kI$`>⷇uV��(� ��]��w/��4�Ҹ$�$��t'8b�~��5����)��8�-���XR���ξ��q�q�,BY`>�ery�%��>B8Ȕ}��y��:�^�j�(��F���A0A ���1���q�D���\�c,��¢^G­x�^�*u�� �<	�wSf�d�
{�Z^ �Խ$?���ֶ�I6Q�K'Z% =�
���wș�{�j��K�� �L�!P�gft�h(���6}�;�����=1쩊
�g�,L�~���]6�Q��6�ZL���}��e�dD�d8�@��a�P��ّ�K$%�G13��{�w��DRŦhHL���B����A������x�v��x������Z�=󗓅�5��bƿ&���}>���k����_��/-�1.j�! =%�s,��`�u���&��nE<P�R���טEC� ��m�}]�"���b��@����j>�L��4wX���Ғ��qdfCQ���j[�x{��<;��o��3tQ�\�%�s�}f �����Xx��޺��z�.m���P=)�����l���	��!������k�T�Kg�^�y���`�r~J:��Y���P)� .��ū�&ng���W>�T��A�@��"C[b�����u���Et�)y��M*Ez���IB��2�+�<֦}Wg
X�����7a9�E�_+b�r��dF�L� 4��="�"�׹�HB�a��n6{Y�l�w�M0:z���/���ȷ�^�x<�U�O��ا���=R�+�I\�	�5�PD����lo��G���wT?&5'�B��y�h.r5Ei�����y
ר��f�:�ll����6�%+~a��M���x�5Mh�ʓ���p�*"NP��oL�;����Zw����PL��o5]0��k��*6-p��8DR�{_���nVEE�9�����|�P�����*�$��- ����q25����F��M�u��F����	9s>���f�{�,��;r5�繚$�/E��+@��kN�΄�}�Ep0�Z�y�L�V��dr��Yi[�)�CÕ��0!kmp��G;��3&�N�¶ۯj��i�uk�;Ѷ4	��s{�����}�=�ɀ®-\�����)jN��<���o��%EQ�����`��-�<u�V{L��V|���'-a�+�*��\�5'��`�-И3�dՙ]}?�+o�3y� ��[��@5��#������4��_v|C��P7�N�Y0=eC��T.u��n�	.b�&h@�5�څ��6���ȓ�S�ߜ�1U��|ݣz٪�Q��=�$������9G��{��*$��Q}-I�ɨ(�W0���O��1��WF1�M��%EK��f�_��E�{�K���j+㆙㫬��M:#uw�dP�����F�a�	`����YH�k#��`�%oΰ��.����:b�aG���;ɬ>+�g��b��Q���D��	����-*"�>[׮'��S�0,f3��51�N&�*;+���Wg����Ye1�X&�T4�iY��ԓ"�|��w0�\k��H��t�@e�M�*C��h���kzQ�Zf) |�Mvl6�h�s�՗��䂸�Uv���}���a���e�}o:T$G* r��) ��f�����[�WhY!�
�����Pi��5:\�j�l�Jѱb(��;0jn_�X-�-X��C��oZoo�(�,�1�[,��>�/���@�h�	 J/3�`!	��^�gjX��=zڪ-x��.�ٙ��D���`��4J��:Z9���3J!��6锼���^g0�!�C5Yhf\��Bd���BrFya�Al;�k+���G��,@x�I"�f]���&�j��\!�6�(Ӑ"�Ǽ���?���~�x�4��.���e�͇�9>X���T�?r6]����թ*����h{���^W}�u���Ao�i���?hP�h�|�����u��8�/z�g�T��-�Xߚ`L&ov�׆�.��	�I��z�n$Zb���E����%P!�)�S�H�J�Z^R�/	 D�`���;/e�l�i�\x�«��$���	/ơ�������/��n������
j*Oxo��G
�7"��:���[��eXh�B����A](z��Y���a)��{&육�{�a�����yos
n�Ⱥ�-B��[g�2x�⥗��Q�ɮ~���f�0�.z_�!���~��U��)WBU��|*'1����o/���4\Y���]��#f6�K���c��=�BJ�hPx��D������F�c0�#��
$�j!�4>��*`1��z�{Ĭ\*�қ�?�he"�fɻ5� Z�@��=Gu}�z�E��{�=�h�m��laFX���戰:AdZ��w�2��>����W�n�_�1�"�$�:?���q��(N`+�%�ض��Vs�4����C���f�I�F�9��u�,"a�y�&�Bhq�9H���:'߅*�z�����(= x�*� � obbs\��/EZf���3��g�}o��?��u�%��ĦM��B%�}bNIW��y�J<�>\�YVË�ݘ����ly���e�8��� t3��4�4�7��4�
O���{*Z�k��۵G4�zA�vǉ�y�� 9͹�F�F���������(#��9�%a��;$����z=F�Fn_8�{�Y��xa��ѝM;���1����iLVo,��E]���M��ⰱ%I�� H>u�0�^��^�(�y��OL���hԙ9����8�WΟz��GM[�*ae��T�����ʪ����#��yBC��:��"��\1+Sr���+q(�C��F��ѭ^���L�I��E�r`p �����:7�c�Y��iQ>�l_��`{5��΢�VL�ؽ�U����~�<�Ƣ������%� b���vfj0�W�Ͱ!�5����If�Fi���(65=k�����X�-/��Æt����X�"���o�Jm+ыm�������R�:al�l���2_ٻ干kF㙘�{N��xJ0�*�'���3gW5SWK��dj�o��zy�-�+��:���t�������eE�أ�d�-�vi�)��ѫk�`Ȝ�� J�����X)��T+�J_��=J���u��i� K��h�*(���7���ɿ�2b�) j��~b�*�>�z�qe۩t꧴t�p����Dp-��p���vRBv��8]C�P#nx�yo��L���YNf������}b�i����� (	�
��^�,a�[��9^�"?7RIi�YS	E��B��'PI�_[D��^W�����X=&´��M �٤�z���Au�h�%��~{�SN���`-����ז%��ݒ�  BL�Ud7H��ջO<IĵN�k��&�����4r}�	�KD�{��m4I�H=�OBQ��1��8�$,���ˢ�	&|6:X�y�dڊ*D#�AҲQ3	qF}S��.�ϖl��hh�>���'��u��8��H��6
?���C�>? ��3�����C=؊�H�IE1��NB	`Tyk�2�Ȝ�D�E({Ҹ
�q��ᙟ��<;H�QlJ�E��x��]�w���Q�[���?�
�򆲙�;d�c����~�s�I�`ӷ�$������|�c���8(�qV�cÏ7��XU�� �r�Z�V��.�!dX�����MC� ���Fo��.�=a�F�u#�r7�\]�@Z�>j��y�#,d�գ���Q���j�B���=8g����R��<�C�g	Is��x�(��Z���	�T��q�>�d}�X����H�1A�e�v�[���E����qN�g��$��={+{�J5��?��@E�Pg�֛=}<®�5��7�a]�oߋKv�ϲ�˴��򅴆����(�����uu�$��?6O:<3��t�%6�S��N�kL���I(LH�B���������zJ��D�q~��U��I��9��=E"�N@n4&��.�։_�&���y�K!��NR�Ps�j���{d8ㅋ x�=���&@ݯ���w� ���i4u��Y�<�"�@?�{7K�OQ�q&��R4�s�����a]O��Q����,ڷv|������,��a�����O��&�iD�;�a {��g{�� ��v�ya�C\�.���~�~�9 &l`2W9�'B��X�}�E�l�1�ys�`�~h�e�P'�	�4�69���`JUb4�8���#�aq��^�=b��C�Լسm�oI�<�uDO�wf\��ӛ�g�o�H��g��ʌ��s��t��8"��?��qҰ�����y��Z?밬�`� ���$��g�����R�?O\��ߩ'�0�"ρ�������.͛Q.1�����%�F���L�zP}��K�]�r����vt�h�^h\d꬚<��	���Hڪ[)�㔋���H"g�B	�R��[�4.�f�<^�6>f���7.<NWG�xN�ja�dc�(�Ϟ9�=��Β���w-���0FĚy�u��!n�yے�H��WHOBh_;���28N>lR�d���Ϋ���6Dm�9$?�V�*!s��G��=9�~���A�\����^�����3ٿ��� �I�*�JǤ���Wɿ���#u!�#�%k��4� o��焆>E���:8W�}�u�:�+�o#GѶ2@���}�@��WD�E���tC�2�b���+�:
�H�פ�kR08P$c�~����
)���	���]�l�#���6_����$�Us,�+�*1l.��%�d2�Zؠ>,�X��U;�C����H��/��h�w�&������?.�Z�s?.������x��Ǆ�����Ǿ��h�;��6F��zp����#G�U��+ U����'��rUL\�M|D��dX��G��=�rZ���F�<���Da�ڏۄ�ƛ&�%a�w�m��<���-�4'3ќI��-|C- ���yb�(�,fb�\�
�����;��	�h��