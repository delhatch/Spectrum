��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k��ib#�Y��&UA��?��?�%|A��͟ĩ�x�Yrl��睇�Z�Ǎ���M+�|҃��4��6��1��O�%����D=�ߝ$�i�b,$��hk��|�FI�w:�
m��:um��q���K4�a��^T�6<�q��2�ŀ$�����:Qy����o���Z��0W��_�V㮽28ߍPU(������$������z5Է�So����{wEr���_��@��G|5m�N>`2"r�'a�'��yF�#�t!N�������S��kb�]��،:��kdX%r��aF��Q`_G!�x���<��u�fo�u��.V��E@#�٣�(�JO��#�����<���2[踾w����h�n�`=�sK�����Y[2��#Im��g�؟a.�S�t��!��ޢR��A��W���!�K�a�]aB4�����_Ut��Q/z���L��;�����M��+/e̗��/-�����Cat��$k�єU��_�z��3?=$�Zt�n$���>�w�E���h؁�@:���r���fў[�%DG7��#�=|L������nT9C䆪�6����=��P*��d���_j�m/Afy�E�~��F���4��N��q�2�r��]��b/j�I��o����9ܔ��s����	4�����J]N򊝳l���\ܘP��!#A{����[سD��\A��Ae|��Lz��|�M��I��ώ�$u�]����"o�:Y�?5�����/G�54U�9J�� �b�dt_������:�H�ʲ�el5i�1~�
�O��}��#�{�1�t���Nc�՚�Vq��}M[^��Knh08�Gp��)�0tP:<ϐ:a24�#KT�h����v��zS� X���n�}�E��~-��%g�  ��Հi6gQ�\��@Ve�k�����\T�#[��\&Ҋ5?t�g0�8�|�5t��:�@g���g�aH)���ך�CYݍ��*�~�J���8WU�+���: �y<�iD��!dX׊�,��v�OX����+�,���0�( Bw�1"P��8�i6=�n6)��F�̜	q%[�P��~n���z�|��7m�a5�ݓ��}����)���iS��R�S���fl����dC�"hDc#�V3G+CZ�����s���#�	r�
�����[Jl��8˲�d�?�8~�$���w�2���uC���As�*�h�'֘�;�?]���Lʗ]�<`�e��\���{y��cti˴��3��KXx\�����e��Qu��͊����/J0nd�t�E�M���J�c�s�[)M߶;JsbR6͌D�l���f�S-��t#9�9�TN��V.���H<�S�8'%�"�Ӝ��Ƨ��D(�(��ΠA�ї�Z�j�A]W��	�vj�@X�uK�c�X�(��@�|6��w�kb��n�f����	��U�	�7/�$Ǫ�2�r��0筸�>��C-ٍ���
�O[ȅG,Sw⟬��3�����[I{V�nh�|³��I������ߺ���z:���j�1H`��G��z�P��f�H����a�Am����1�͠5O�~��60��Z}� a�Wǚ-̠��Flb"��Ԅu���	ЛQ�a<?>��3��W�����Z@1\��Ɵ!�+6c���P�g0��_5�8,!�᧖H��3$�Mq��-+�v0�W��������m�e�AZ�b{0�g��+�_�*km���2��ţ�>4�
5ϒ� �"�S��ɛN4��Mr���$� :yH���&5s"L�M�uD"M�HR-�����~���V�e_��O��꡵��oA�ۮKQ����x��Kh���]ġk���2�Ψ�C[g7LZb睶G� )��Q���� ��ª�>e���,/�%�3����z�D�cc!�j	��>[H���I�4��M,��#�ݏ���(F�ȾV�+�eŗ3���'�7�����p̮IE��S0i�Pu�a�RR� �?Θ�#�!�3ا�5?L��W`���i��+s����u�hb�f��gi��G7�)�9���ifyw�$����;�˷�A7�Քz��+k��~��7ab3�����vf�d�{E,��c8`jnm����?�d�@a]�mF���oK��<r@Mg���L�;=��jP{�"���B4.�?2��=�A�&�Q��9\wlj�d��`�r�H�㑛�¡j�4��Q� E7�t�2,���9O��(�/�9\~���@���Q4�����ů�1�;F�xf�t�o� �Ρ�1"|����7��!B�v�i�h'}��KD7
#|ʺ��6)g�M�Ŷ�K6}�� � ��dE{���/���q�V��ך�o�@M�'�u]=Q���� x�|	߮n�ual�Ƿ��{LG��%!oL̮V��u��e�F�t>^���6N�q�N%�҇�,0)�Y
G+%�������2�J?�2��D͗li[���3B2��=yg�M�͌&���-�0~tE��i��&8��!�L�ǤΩGĔ�X[�0$�Z����7R�M� r}��({F�Y+�.������n����������1v8V.�(�7��;�}�	~)���@�ȿo��!� �}).k�!������9��=���`��ow?�����~_�Tޮ1�U`O�(���L>��u��d�9m=rSD�n�4����\V�"j�/A�J�uX����T}�|pFwg|5[��XZڬ�اw�D|�C�t�2�s$o�V�Hbf���㽥��:i$mט�E��DWg�<H�����~�{�;�H5dpt���p�ǫ䭊�q��YS�_>��X��7�{ir�\! ~A�zU�t>G��R�KO�������4Ay�/�s�7��;�נ%�tp0~!l������k�ZGI�ߊ[Ro+|�C��ؙ-�_���(��K~��?T������B�vpJ�j���iDSޖ[�����V���"N�ёYW������[k"prZL��Oel�a��"&/7M��%�� p��i��A7)��	���u��XבN<�I�������M�.bAe��Xm|�.L�ΓW��U�lyTBl�8i�,�`������LI�vЅ�E|���C��  mu{��j�Z�:?,�u��aa7p�M�S>Ǎ@�1��5Y��=���H�Ȧ�bW������L��'�&��K���n���=��FB�E�4�(�x�̓��M�a�QU4BP�XRE�w' �5U��ZT��5�5���n�	90{�(ǒL�L�VS7j�),c?��30zdH��
���e�+*aD�E���<}��^��GJ�$��h����`d�!�	��h�R��J�UWn*�����ٵ�������XM��+��L|��̔h|�y-�%&�g��#�����u1�tbI(�%>��00�~��c�6�ʳ�\��f⩓e�'�	$�'ɂE��&26ߔ�MEDO4�w0��ë�~y��XtA�̌��6�sR�ڲ�>S߭5q�N,�'N�`�
��G���9��u��߸uR@q܊vn�#�,N�F����.��^Z!O5̌~B��4zd��`M��{�@�F����5��s�s��V��jyT�e��{��Em�xv���IJ��Q	B����]"z[:��v���ʡ�r�m��v�_) x���������3�)�%����W� 42Ȗ��F��ǝRUC�O�J,TE$�x��~��Ϋc�};�t�,{Xl3~A=#w�A�^_��o��-U>�d��P*}��t�r�?��Ԉ��1rA�.�(e��
\�(�t�T��r���"�*;�G�`�aftT�B<���V�1pb����x4�3%*�����
��D�L+�6{���.[J�5��ȥ֣ao�.sf�z��`�e�h[�L��=���I���Trs���|�z���%f2-�Ǹ4}جgj\�PS���w<(h�Â'���1��ri$�7��L�����e��1h�t+@)r�
v=L=�oZ�F4�
2�	�<M�3;�Y��]6˽[��:KdBc��	Y���w�^~߈˼��~�=fT������Aa��,tx�4(;s{a�ԓ��U��G��NH���S�$4!�70p�o,��
Rѐ���o9�uQQD���s=��Y�� �_�*=�?uy�4�����n�y5���~��p������g��Ĝ�%�ӯ���M�]_	fB�Y��>�>�p5�'	k�w�.����H��F5B*���
&P�r#��i鉍�u�tf��K�0o;jDx���rW ���i��@�еߧ����V��r�։����{�1Hs� ����]��F��	��o��q��=<#�W�9����.�v��W��wH	'Ѣ	'�����Z`�5&%�?���`BS<�r���,;Ӡ�"�����`��AL��8X�Ӫ��]�!�+rㅬȻ��h*<;����8�xSu8�����#��)�S�G���Y���	���x���c��1��>�҈��7��og�^�P�$-�Á��F��9R1�ĆF�a9P��LP���j�Q�z`�[����]}&{j�^��<)|��sa	��) ���(V �Ճ�CQ��.nY@I*ܣ�����
�9�-�QG@_���}9�z�٫���U��c�	+}�=hY}@�T�>���6	�#�|J�!������,��
��16�/cN��nrD�8�ӑ�WU�\�]���=�f[M�⿢t�To%���Mi�	I�y���s���q��t���O�f<ys[�C&$�Knڙȝ2b��tY��r_��=��
���M�6����M�W�Z��"A�ݟ����	�6Q�l�Id���[|F�]U���hu�D��\"�I��ۈ b���������bvM����q��	��J�$j���a�B3I�3�1�O�Ma\�Y�Ջ�3O|��l���zGd3���*���Y*N�v�0���}�!O�15{JDr��W
p�u������}�EP��}��E�yBc���<�M^u��iK�n��_}���|<�/~�S�/��q! kg���Eec��(�BC*d<���9ő׼�!(Ⱥ�H#��͋�.l�[@&|"A�?I��S�� gcBPKW�V'S Y,�c�+1�;�mv�����IػV}k(���X���VjD��Gmm�