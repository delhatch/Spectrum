��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�Xuѳ����\�{J/�(b4&��kxBa��(q�_�p��f��*�>���Ù���2�0��y�/���ͤ��������z�T`kc9��N��'�y�`�P<d�,bL��}������ך�]PV�����Dx|�|	}�#Ƙ������ ��Q���z"E��V�&5���f�(�f���ŗ��o��f2�}�q�e�Э��א	��*��9����G�̔5?���&Ϭ���x�\�>�����M���OM׃Ad��=9��o�1	���]XEo��|`�о���7�p+�JN�)�~ZbM�(qЩ&+�=��%�W��б�i;NЃ���q�wK�w�܊U=�%{�š������y�(p�1(F&˂�v=���I�8	1���Ņ�����>�ͻq@f��z�;���#��A���^�X�w���߳P��|�/A���"��4����1�s�E��S��"N��������Jw�in�i��\��3�Y_�`�X'_�Ku~W[J�����d+Q�-�K�g�J7���0��ܴ��?0.��@G�`o��i�C$C��H�SJƞ�J6fm���]Ֆ(�%��T�3�^�+���R�䭤��fK���wc'sfp��V�#6��ݜ��L�xTO�Z�������.��#ך9������i�\�1��Ά��[�s��0,����^����S�!z�m�Ƴz� ��1jgH�wr��^MZ���~�U�����R7m��B�1�W=��ָ��Ep��+�6 A��U!����G�<�k����i*����^�����RE�6v��(�zg`!���ay������?ejY{��B�<�ߓC�5�EA�v�4��`^��7}.�� >9���k]]�h�H�8���n����L�b��������S��W#�`�Q�mP�5��f�[.�� �VP��=p��	nJ-ͫ��"o�F��4��� �������p
�X����q���x��,����
��G؃����h�6�0��"O��.K6X/ #􌃡(�����:�4N�����������l-��������`讝.��c����0�~\���`Cʓ�S����EL�y�l�.c&M�M,
0�w�ѧ��m�����5i��=GBY{ �(>�d;
{!t�6�k���]�+%fs��������o�h�����q�����#ˁRVPʁ�!�(�� .r��s'�H�cd,��� �WKw��R
*����Ԉ%Nt�� =�<\���z�Ԕ�rϐC�.57-ג�erW?m��\d��Z�}�S�R��O�u?����N�ln.��jU�2��j��1շ��aV�\_��n
p�&~�Ȭ���r��[Y٣[cw2�����@��7b�j��71���"�%Z�����8_���$��{���(9z�����Z�y�Z]ZķZ�f�����r��k��	�U��z5�*�ZŢ�1:��2|���s�=���|��w�S��6F�<.z�����;֘�<�ASx�~�����	�00к\���:�xs���v{���41��o�R���:��u�GHGs�(�2��S��W�Qg��>E���3yQ�:b\�U�����V�J��u����c�,�1zHܑ��(:!<�Z�O���Ki���V�uh���b�Q�N���|ln)���v�}�i6����A�1԰,�� �^�C�e]=�	pf�Օ�z�V 4x�L�6�-)�mdC���g����e4
l!�P���SG�4��rxs
��!��Ԣa/��~�&4ϣj;5U�݉�]��E7��k��CXd�z��������� �m
�r�X�=�a�C�{_��X�)�ҟrL�a>{	����ܖ�HU_%�."Bu�b��-	��a�J��M)"�8��� �T���|����1��n����1�5��W"�w'��G&�a9�<�TX�Ζ~�	�k�1)&��ީ�O_Sl�a��/�d��O�x���Ӄ$�mH��'�����ƾ�j#�cU���vț��m %�,g$E���8��'�IE�^�'K;A�LD�|ҧAo�w�S�f#I"�I�л�zwZ�~֟�r���QF�
�/,�B6A�޳fѩ�2��Q��캆���"��Q���:W�00�"�F:< ��27K9}���0T͔���h�,oL��?0(|���Zt��'l�h���2O�t��I)����-����Ol�s�*#f�ˌ�̖�M�ޜb߸�����]M�� ��T{���,��|�����r%�nz���0m��?��X0�D��I�?���y��ʩ�\��ٯ�D�<lnOM�k-e��5����Tʹt����h���xHT?�FxK���l;ޒ���#�w4�=g�XF$#E���ϱ���SZ�q�֡BF����XwG���FDj� ��� C�Z�{���f�S��tZ�.��k���j�ṧ3��wLF�\�?SJ9����`��m��h��X��C�i���l�0���@V!i|�=�e����B{�p�-�\�m���7/�tq,��q��K�ĎXi��LE�-�[��g����fj~�xܣP�4����!C�r��p��!�nǨ4���ȹG��fG��{$���eRA���ښ�2r���� ;P�~����.�����N~ �u��I*`O��s����~��,F9�"!懜]�O�S0#���XE�OK�fZ4� &�d�A$����o�J�� K,��:8�8��Ů~��)��q����F�A`�����l�y�S`�J�����G�M��X���L���v
�RI4�P`�q��^�6�t�̝t�&�|��5�_���k`�#9���4�s���k�p�� ,̗O�F���x�kD��&a.�T9�3-�L����.��C$F�S��E�7�@���ѭ��C��Y���铸t�;�!���C }pVY��ī^����WE�xnWh��-0�uv�GB�O
-�?�&y�NΆ�
��(&h0N8�$�v� $�e@O�������]*��q]��_2� �ub���C��~��C���1[�	t��~=��(>\
���lC425x7�?��1�~�;(�@V�
��Fջ�vu�����v��Uq���8�Yx�u��FN5�P΂��YOyq���SS� �qZ�R��$7�e(XW(���tˎvǃ�2��3��pѭփ]���$)�T?��6絣l˓�2���4��ؗ�����*ϒy�U�1�[�*[o��2��I��5��q��N�|�Mgk�3�0��(s�B�>�	��/8��aB)���z`�Kj"s,f�1+zSD�m���K��4@�����ˢ����5�� ݔ��ݷ����\����Р�"r�O�������:�Q�"T�*�0�����,��b5r�Ĕ"���|f�,�r��ELO����mM�O�4�n}�c%�&#g�&��x���YX�"%5�]�P^���F���'���~n�o��@	��m�9�r�_�YLKx|��_��ݼ�����ᤂ@� �j�%7�r��� Q�3+RR�'5����jDK�?]�y�Y|7*���ڏ�d�HE+���S����R��<�P��r����X�\Phׂ�0'�@�&��U8}��Ǌ��#z���1��l�;TJ>��?�j`a/zQ��`���K�	�C }�$dC�s �+q(��w{�هx{����2�g��9�^�]#Z����q��$�"��HR��Ŷ�*��x��`�+u!rCGk{�J��Lدtz�8���@73�� 4��
�&?T��^5~F�	S�F@����-�hfO���ʆpf^!�ʌ��~��\0{=]CŐ�f�����5�zL�ax�)K�F�J`8��Q�%�3���g���<�����.`���P��Z���Q^FҮ�Wp��s��8�Ax��N�鬠��(�J��.�� d`Ò�V@��#�:Ӷ8�� G�.��TI~�Vy�b�&�~2��:-��˧� HP'7�����Gz�漑-IߧԴO���Sgf"�����LL��z��������=��9T�ܷ�U����r��%�e����Uل_�R+�"�ŷ�I�{�PV��a��7��R�i���4�������
.�j�GZ���c,JNQ���8e֧P�Q��� ����%��l'S�ށ�����7�dR�%����mo��4~���!w4�\�~4���|H���ܓ[36/�'� �� �%XS��_��+O�Hceû*G�ám8W)�Q�{�(m���;��(�G~ՠo���
�����n���sV�����H^��Fu����N��J�ZI�/>"]!	\���#00�W]aA)� �gZ�4;m�l����k������� p�?|8�n\W%"- q���r��iǭۚsj���e��<�\k=� +���W�<o#��[��yvɏe��s�孛�X��)[�|��Y>�rm.U�~�f(Qȸ�T�#�aàK��6�����Ǟ$u�������`g=/g^y�w�-髻�Gۚ=��m`-J�Ý���RuS����]fO_
B�\����22�m]����k���f4��q�<�[ ��1Zi�.��~A�?!�K/�u�]=��!cƊjS״}11@ml�Ï��XSHF��jX��kI�O��`�2���*�Ѱz���W�.�.��������rf��zN�e2��˄~>
� Ĵ��X��:��\�&c���.�i/k5d�I(�	�#4�GHǹ��+ud�c8�]�L��muE�Uv��Т��a��|k8�-K�������S��V�rG�砼���v�:��������c2��C.���^=�4���«� ��r��V_a��a��4牕�V��#��Ef��?��[=���x���4��K�F�I�R��76�f��g�%�U��1��Xh�a�[�"��s.Օ�kǩ��f�ehɍ �si����:�E@.\��L S��S��J6��je۔'x�R��	�����Oo�e���h���{ :t��u����m�K��v�~���[|���Uk7��;����MB��t�`1�:V��[x^+ע�-{|'�?x?��/<hǚ�$z�4�ql��:(zQ�D����c�1�6��&2ޮ]@ ��%��Y4��c���͘aC�q�S�{|���u3�����8��� #��l�>���m�ah�()�O(v��� ���`�-�]��]�&���xd(07��a�Vj1R�+��Z��b��Y���t���*Di�o�w�<Z�Kr[�,;�"t��qB�c5��q�V%�)S�]��Ro5!-����g�v��BP�_��Y^J�&�A����o������g�I���{�������T�kV��0��?�
7�Qv��"çxʙ��(�J[�N�W�,�O��c�pi����������FϜ�l�@��ò
�.vޓ�Fˈ�r��*��m����d���M��a����_C��"���q݇��s(���Z=�+$tv�+�r��>��Nz˷-�/�wb�e:i|D���i�8�t�gm��?�64W���@����X���V��R�K>&a����27��j!<3s���&�:!�Nb<�F�Ӈ��$to}��ח��V�{�g��cC'~X�.ntxx��@����F��d�j����H����O^Y����滝H�����y�6��PEo��T	'�A�>Bϗ6۽6%���~��0C�jB�/9��E���B_'�bxJj��Q���u��H�'� �W��1o��u9��+������ʪO1�s]����p����@n�fk��"�p�2 ��C��u�c�W�|��{^�Xju�ϸ <Uv��\��%i�g^�����6I��<_:��;��{(4��C��t�L��;9&#�(��k����saIv!��U&��&� Q$3�8���Ձ���g4be�D
�^�I+��0K#.�f�U�z�?Z�b�ތi�!/�}��k�)�`3^R�UQ{���~zm_&igXF�o]��To���ll��#��p�&_-��3W8��Ð�L�R�I@�^�UUl���=Y�k��gh�����{ERz4k���M�
�@\���F�����nI}� ���	�U����E/.��T����n�<�u�;mp7����oEI�tA{5%d	ēO�l'�_3�Ƌ�_���^��h���������gsS���pO�;���%�+���.+Z��3*���A�Ëv�	b��(��\�������Y�G5�IVӹY�9�n���6>KQ37^T���i$Ѱ6=�h�Ptx�O����"�U|��&G�Õ���p���Z?�.j+V�^q��r���6��!�IK!;xg��DHT���Hp��b����0<�닳g�y%7�(����=Mj�IQ���{�b@	c��:5?4O��ԏ#���HC2��Ǔ�ϕ�"��`�Fb������}��Og/�(#C$:%,��կ��2�L��z�xm��1��d�`ˍ<���?�Vf�����1<���T�O��YDG�*�؄�Oc�-�fM�i����5�k��xG�� ��7_��\F��q!�g["����:܂��2�5�c&�\dv�ym=��}a��B ~r�)Ɇ�N�N�%ڼ�v�xt��#��BaS[g��d[v>�Z�������.G����?�X��c��cM���N�$B�G�@�Eo�"��d��G%	���tW�l�O=Nq�޶P �q�����E��������^�)�� �oMG�B���#�D���\g�3�+�����~�/Tj\���|�ò���
ze%��#\�g�����Rc���Բ Eo�
��
�D����,v�"C�m˙Ԋ���h&��M�\ng���㛎��Z��D��i�������h��Xļx�} �c�Ȑ�'�a���R�\Ql�5o���;�U������;6���`��G����3߰�m���_� �� G��S���`���Ub8���EiWsw���w|;�mKSK<-��z,�Q������H�hA�R)H~B��0Tn�"� �0 ���2���)�^���|H���W�&'{�u���Ï�^��;��Z�1�]J�Z\���9��p����6��|� ��)t��	����0K4�(�R�8�K��K��{�Ō�&�P,U*>-����%:�萏��?������)�+��v<# ��A-�N��o�`�S:0�"�b������3xK~X��`�U�r>1�����x ��3a9�����|J3����E�ְ �kn��{b��5�F�q�����>I�I��$��7��0z�������l�W꠨^�%tm�V��h�5��n�(n��yJ2�	r��ȯ����@�l��jm�|��8O�e��Xk�}
o��Iv�iYA�x�s.�p�aĢH�K&#��Q��\]��^�m�Y5��g�?u��۟m�����,�6,y�	w:mF��u����+�n�k<l�2���!�K!��Lb��7LX������s��V�^��9\*��T��L@�$�T4Qj�V������52$d7��dc#I Փ��$�(ݙ�$�v��Z9'D���̦:����ysǴ�m6��nH�/\Ð��m�<�	�Pr�_���tDzl��s����r�^݄��% v[ׁP@�0	S���w�C�)	�����wz���'�D.C*{���w��Lx���+�*Y��I&ͮ�D\�L!y.D)�.F��UKMi��zhNi�9e 2S�G�9��C�EN���yQ��e_���Y;� 3ۑΙy�	��afo�Y�V���хQ�KP>�dI�7Z6��#fj��f���X:��+���r�����d%>Ϧ�5��M��AA�$�����ZqB4Rф�a����<�����`�����w42T��=�vQ��1o&���O"�C�\�)�to!C~x�f�,2��n��@�cf��֬���m���M�T�O���P�s��|f��0\���,��h�@�?1̕Q�8,>�Ξ���)w�gWږ����ߙ�i �h�͌���$�{ɒI�>��?��a��^ծO#U	brgrb��P:��|��y�+,."Х� �H�A*�q�1���
�~Ӎ������߀�]���TM�9��= �ן0W��&y�����,�0��vd�f�=�;B�^ �j1���5H'���(AL*��Թ� |i�"0�����O���A(�r���f��	Vw��P��[~�!��v�-���띣��^�9���>�H��
�4��`��Qb�w��_��
��?��DK�Iʌ�W@��E��Y@
#�w�k
<����pAm$.
���R��ҡ�U��I��Sq��-������
���s�Q�*0إ=oܛ�����b�N���+$g����;�ߴ�A�g��4R������M������xÉ��{������`Gs�~�����k�e���p�険2�)����h9盧�]������ђA�����w�!���������%��6!���P�����t���̬�t�s��	a�\ȇn�斈�� �q�a8��'Ŏ�F��(��r!���Jxr\��Zʾ�1'J�:M��}g=�w�F]>i����g�@���n�g�Ū����Ew(�mH�I�w���A�P5k��*�3w��Pn9	\�}�I(���;t��G���r2��=e�a8�?Nu��d��A�.8W�ʄ<�|'��$Ѷ��1k`*��"�.��Qg7��5��}��ίL̾�Ų��h�z�3,z.:�9D|��B*=��D�PtM��^;�����V��O�؀�P-DZYeč��P�/�v�w�� �h���J���AB8Bw��9�g��Q&N)�m�����"������7�$�rx�<�F�^a>]��G��K� ��1��װ0S�L`��P��IP�,�ep�k@6�-���b�&BZ#^�3VT���Xk�ZI�Y�(#��w��meZ�^��{:1c�vi�p�uq��?����t��R���6�ƨ��Y��c[s��s���C�֢"A(:=�⟧3H��&�"�Aߠ"0�C`��)e�D�NfY��#�p��LC��[c�!�����8�)�ȟ����L�i�L@�̂(��N�CF�~͑��� �4�iA���6Nw��y��e+ZL��:獭 ��E0z<�jK���k�pX�H�{� �"c��#V�خɁ�tXL&*td컀�xY�}̈́��*�%��>�;@	A������A70���~��#Y�Aw�����g���U�����T���-e�h���un`�W��#���%1�3�3����8�)Tj"�Up1���&\&��u�uQ'��E�+Ss);�'q ���� �
Țƚ��/�"��j�r�&ܢۼYαk��C-��� ���r}��ψ��'��	�s18�ST5�]<>o����'&�E�x����#�5�n�H�)�R�8WgP��y7hf��|mn�V@��������+��p2�����#E:��'v�Lf�x^�<k�E�.0"�g�0�`<�DU�4��l�uL�N�����Kf����Ocd��8i˚��U���T�9�D9w�	M���ſ>oWl]^SӲ%�%�8�k%5�
]5D�xHH�6�[����f�P��$h�Ec�����3�WL���,�ŭ����#S��9{���;�p�����y@AK�{)'�~�Z &�6�5������.�8/Y�>s�zs��f=�����`���+��Q�w��n�Z�Yp\��˿Hube��U����w׀�����[y���R��S���y}Y�:�QG��Fb��rO+/�e<��*��Cm��!)<�\�*%3K��⣪����D7����*ي�"�]{%ݫ�psގ6Y����+ �pD�v��F�h�M�����]�����o�#�l��E\|"w,��[�
�>�~��!������Yi���� �y}X��T��T��D�Q��TϮٓ���0��>ՙ���iEd:���O���H�D�j��H�����K� uffV-�@�s�O7�>�D�&��z�8�6�zf;�b��OZ�ڑQ�yF�p�[�n�O��>_@?��E�&0|E�S�܎�}��E����u$��	34w�0�3�9�Bw$��.��r���[���W���<��Yͦ�n�h"��F���˃��ZE���� 9�5��Y��J˖|a��)�[
"����X�t��i��ѷ������{�z�Э��H�2��L�3D�@+���M�\:V�Q
�A��֠���U���Bp��K�V[:M��0���:罍TVH�(
X;B^]�Ezq�:#Fg��冲�۸k��ˢ��'x���c�hI��9,���aB���s���T7m��J�6iE�'��ɱ���ͦ)G����
�� [ \�U5{�cb��́訓�DP���T@�,O�� �Ǆ_��<1�u��[��,�q0�ɉT�/ �B�đb/c=�M�@TryC1�[cm_�F��K"�@���x��a���{�r�v����2� D�u#2���;�������/��0�'�ߦn���K��_,W���fx0��#e�Y��K��1��=�U��k���)e]��5���f��g��t�Z(��A_aj����4Y�{�i��e���̶QҪ���Rl���	�<)71�0�(g��2����1�B,QݒմFsh�W��Ď�NҒE�`�~e�6�(�^�a��r�,!E�*������ ŬJ�zj0ͳM����'#y��Kݣ3��%��Yp4:N �[�g�_*��J�N�0�8���?