module Spectrum(

	//////// CLOCK //////////
	CLOCK_50,
   CLOCK2_50,
   CLOCK3_50,
	ENETCLK_25,

	//////// KEY //////////
	KEY,

	//////// SW //////////
	SW,

	//////// LCD //////////
	LCD_BLON,
	LCD_DATA,
	LCD_EN,
	LCD_ON,
	LCD_RS,
	LCD_RW,

	//////// RS232 //////////
	UART_CTS,
	UART_RTS,
	UART_RXD,
	UART_TXD,

	//////// PS2 //////////
	PS2_CLK,
	PS2_DAT,
	PS2_CLK2,
	PS2_DAT2,

	//////// SDCARD //////////
	SD_CLK,
	SD_CMD,
	SD_DAT,
	SD_WP_N,

	//////// VGA //////////
	VGA_B,
	VGA_BLANK_N,
	VGA_CLK,
	VGA_G,
	VGA_HS,
	VGA_R,
	VGA_SYNC_N,
	VGA_VS,

	//////// Audio //////////
	AUD_ADCDAT,
	AUD_ADCLRCK,
	AUD_BCLK,
	AUD_DACDAT,
	AUD_DACLRCK,
	AUD_XCK,

	//////// I2C for EEPROM //////////
	EEP_I2C_SCLK,
	EEP_I2C_SDAT,

	//////// I2C for Audio and Tv-Decode //////////
	I2C_SCLK,
	I2C_SDAT,

	//////// TV Decoder //////////
	TD_CLK27,
	TD_DATA,
	TD_HS,
	TD_RESET_N,
	TD_VS,

   /////// USB OTG controller
   OTG_DATA,
   OTG_ADDR,
   OTG_CS_N,
   OTG_WR_N,
   OTG_RD_N,
   OTG_INT,
   OTG_RST_N,
	 
	//////// IR Receiver //////////
	IRDA_RXD,

	//////// SDRAM //////////
	DRAM_ADDR,
	DRAM_BA,
	DRAM_CAS_N,
	DRAM_CKE,
	DRAM_CLK,
	DRAM_CS_N,
	DRAM_DQ,
	DRAM_DQM,
	DRAM_RAS_N,
	DRAM_WE_N,

	//////// SRAM //////////
	SRAM_ADDR,
	SRAM_CE_N,
	SRAM_DQ,
	SRAM_LB_N,
	SRAM_OE_N,
	SRAM_UB_N,
	SRAM_WE_N,

	//////// Flash //////////
	FL_ADDR,
	FL_CE_N,
	FL_DQ,
	FL_OE_N,
	FL_RST_N,
	FL_RY,
	FL_WE_N,
	FL_WP_N,

	//////// GPIO //////////
	GPIO,

	//////// HSMC (LVDS) //////////
//	HSMC_CLKIN_N1,
//	HSMC_CLKIN_N2,
	HSMC_CLKIN_P1,
	HSMC_CLKIN_P2,
	HSMC_CLKIN0,
//	HSMC_CLKOUT_N1,
//	HSMC_CLKOUT_N2,
	HSMC_CLKOUT_P1,
	HSMC_CLKOUT_P2,
	HSMC_CLKOUT0,
	HSMC_D,
//	HSMC_RX_D_N,
	HSMC_RX_D_P,
//	HSMC_TX_D_N,
	HSMC_TX_D_P,
    //////// EXTEND IO //////////
    EX_IO	
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input		          		   CLOCK_50;
input		          		   CLOCK2_50;
input		          		   CLOCK3_50;
input		          		   ENETCLK_25;

//////////// KEY //////////
input		       [3:0]		KEY;

//////////// SW //////////
input		      [17:0]		SW;

//////////// LCD //////////
output		          		LCD_BLON;
inout		       [7:0]		LCD_DATA;
output		          		LCD_EN;
output		          		LCD_ON;
output		          		LCD_RS;
output		          		LCD_RW;

//////////// RS232 //////////
output		          		UART_CTS;
input		          	   	UART_RTS;
input		          		   UART_RXD;
output		          		UART_TXD;

//////////// PS2 //////////
inout		          		   PS2_CLK;
inout		          		   PS2_DAT;
inout		          		   PS2_CLK2;
inout		          		   PS2_DAT2;

//////////// SDCARD //////////
output		          		SD_CLK;
inout		          	    	SD_CMD;
inout		       [3:0]		SD_DAT;
input		          	   	SD_WP_N;

//////////// VGA //////////
output		     [7:0]		VGA_B;
output		          		VGA_BLANK_N;
output		          		VGA_CLK;
output		     [7:0]		VGA_G;
output		          		VGA_HS;
output		     [7:0]		VGA_R;
output		          		VGA_SYNC_N;
output		          		VGA_VS;

//////////// Audio //////////
input		          	   	AUD_ADCDAT;
inout		          		   AUD_ADCLRCK;
inout		          		   AUD_BCLK;
output		          		AUD_DACDAT;
inout		          		   AUD_DACLRCK;
output		          		AUD_XCK;

//////////// I2C for EEPROM //////////
output		          		EEP_I2C_SCLK;
inout		          	   	EEP_I2C_SDAT;

//////////// I2C for Audio and Tv-Decode //////////
output		          		I2C_SCLK;
inout		          		   I2C_SDAT;

//////////// TV Decoder 1 //////////
input		          	   	TD_CLK27;
input		     [7:0]		   TD_DATA;
input		          		   TD_HS;
output		          		TD_RESET_N;
input		          	    	TD_VS;


//////////// USB OTG controller //////////
inout           [15:0]     OTG_DATA;
output          [1:0]      OTG_ADDR;
output                     OTG_CS_N;
output                     OTG_WR_N;
output                     OTG_RD_N;
input            		      OTG_INT;
output                     OTG_RST_N;


//////////// IR Receiver //////////
input		          		   IRDA_RXD;

//////////// SDRAM //////////
output		    [12:0]		DRAM_ADDR;
output		    [1:0]		DRAM_BA;
output		          		DRAM_CAS_N;
output		          		DRAM_CKE;
output		          		DRAM_CLK;
output		          		DRAM_CS_N;
inout		      [31:0]		DRAM_DQ;
output		    [3:0]		DRAM_DQM;
output		          		DRAM_RAS_N;
output		          		DRAM_WE_N;

//////////// SRAM //////////
output		    [19:0]		SRAM_ADDR;
output		          		SRAM_CE_N;
inout		      [15:0]		SRAM_DQ;
output		          		SRAM_LB_N;
output		          		SRAM_OE_N;
output		          		SRAM_UB_N;
output		          		SRAM_WE_N;

//////////// Flash //////////
output		   [22:0]		FL_ADDR;
output		          		FL_CE_N;
inout		       [7:0]		FL_DQ;
output		          		FL_OE_N;
output		          		FL_RST_N;
input		          	   	FL_RY;
output		          		FL_WE_N;
output		          		FL_WP_N;

//////////// GPIO //////////
output 		      [35:0]		GPIO;

//////////// HSMC (LVDS) //////////

//input		          		HSMC_CLKIN_N1;
//input		          		HSMC_CLKIN_N2;
input		          	   	HSMC_CLKIN_P1;
input		          	   	HSMC_CLKIN_P2;
input		          		   HSMC_CLKIN0;
//output		          		HSMC_CLKOUT_N1;
//output		          		HSMC_CLKOUT_N2;
output		          		HSMC_CLKOUT_P1;
output		          		HSMC_CLKOUT_P2;
output		          		HSMC_CLKOUT0;
inout		        [3:0]		HSMC_D;
//input		    [16:0]		HSMC_RX_D_N;
input		       [16:0]		HSMC_RX_D_P;
//output		    [16:0]		HSMC_TX_D_N;
output		    [16:0]		HSMC_TX_D_P;

//////// EXTEND IO //////////
inout		       [6:0]		EX_IO;

//=======================================================
//  REG/WIRE declarations
//=======================================================
//seg
wire        HEX0P;
wire        HEX1P;
wire        HEX2P;
wire        HEX3P;
wire        HEX4P;
wire        HEX5P;
wire        HEX6P;
wire        HEX7P;
//vga
wire        clk_25;
wire  [9:0] vga_r10;
wire  [9:0] vga_g10;
wire  [9:0] vga_b10;

wire        reset_n; //reset

wire clk2fft; // carries the 10 MHz clock from the pll at this level, to the fft in Coproc_Top.v

wire [9:0] mygpio;
assign GPIO[9:0] = mygpio[9:0];
//=======================================================
//  ARITECTURE declarations
//=======================================================

assign reset_n = 1'b1;
assign VGA_R = vga_r10[9:2];
assign VGA_G = vga_g10[9:2];
assign VGA_B = vga_b10[9:2];

DE2_115_SOPC DE2_115_SOPC_inst(
                      // 1) global signals:
                       .clk_50(CLOCK_50),
                       .reset_n( KEY[0] ),   // KEY[0] is a pushbutton that is normally low
                       .altpll_25(clk_25),
                       .altpll_io(),
                       .altpll_sdram(DRAM_CLK),
                       .altpll_sys(),
             // audio signals into the system.
             .audio_global_signals_export_adcdata( AUD_ADCDAT ),
		       .audio_global_signals_export_adclrc( AUD_ADCLRCK ),
		       .audio_global_signals_export_bclk( AUD_BCLK ),
             
             // debug signal bus.
             .audio_global_signals_export_debug( mygpio ),
             
             // clock for the FFT portion. Not sure how fast this can run. 10 MHz good trade-off.
		       .audio_global_signals_export_fft_clk( clk2fft ),
          
                      // the_key
                      // .in_port_to_the_key(KEY),

                      // the_lcd
                       .LCD_E_from_the_lcd(LCD_EN),
                       .LCD_RS_from_the_lcd(LCD_RS),
                       .LCD_RW_from_the_lcd(LCD_RW),
                       .LCD_data_to_and_from_the_lcd(LCD_DATA),
                        
                      // the_sdram
                       .zs_addr_from_the_sdram(DRAM_ADDR),
                       .zs_ba_from_the_sdram(DRAM_BA),
                       .zs_cas_n_from_the_sdram(DRAM_CAS_N),
                       .zs_cke_from_the_sdram(DRAM_CKE),
                       .zs_cs_n_from_the_sdram(DRAM_CS_N),
                       .zs_dq_to_and_from_the_sdram(DRAM_DQ),
                       .zs_dqm_from_the_sdram(DRAM_DQM),
                       .zs_ras_n_from_the_sdram(DRAM_RAS_N),
                       .zs_we_n_from_the_sdram(DRAM_WE_N),
                       
                       // the_sram
                       .SRAM_ADDR_from_the_sram(SRAM_ADDR),
                       .SRAM_CE_n_from_the_sram(SRAM_CE_N),
                       .SRAM_DQ_to_and_from_the_sram(SRAM_DQ),
                       .SRAM_LB_n_from_the_sram(SRAM_LB_N),
                       .SRAM_OE_n_from_the_sram(SRAM_OE_N),
                       .SRAM_UB_n_from_the_sram(SRAM_UB_N),
                       .SRAM_WE_n_from_the_sram(SRAM_WE_N),
                       
                      // the_sw
                      // .in_port_to_the_sw(SW),
 			
                      //VGA
					        .avs_s1_export_VGA_BLANK_from_the_vpg(VGA_BLANK_N),
					        .avs_s1_export_VGA_B_from_the_vpg(vga_b10),
					        .avs_s1_export_VGA_CLK_from_the_vpg(VGA_CLK),
					        .avs_s1_export_VGA_G_from_the_vpg(vga_g10),
					        .avs_s1_export_VGA_HS_from_the_vpg(VGA_HS),
					        .avs_s1_export_VGA_R_from_the_vpg(vga_r10),
					        .avs_s1_export_VGA_SYNC_from_the_vpg(VGA_SYNC_N),
					        .avs_s1_export_VGA_VS_from_the_vpg(VGA_VS),
					        .avs_s1_export_iCLK_25_to_the_vpg(clk_25)
                    );
             
// Configure the audio codec on power-up/reset.
config_codec codec (
   .clk( CLOCK_50 ),    // 50 MHz.
   .reset( ~KEY[0] ),   // KEY[0] is a pushbutton that is normally low
   .i2c_data( I2C_SDAT ),
   .i2c_clk( I2C_SCLK ),
   .xck( AUD_XCK )    // becomes "AUD_XCK", tied to pin E1.
);

fftpll thispll(
   .inclk0( CLOCK_50 ),
   .c0( clk2fft )
);

// Tie audio input to audio output, for monitoring proper operation of codec.
assign AUD_DACDAT = AUD_ADCDAT;
assign AUD_DACLRCK = AUD_ADCLRCK;

// Flash Config
assign	FL_RST_N = reset_n;
assign	FL_WP_N = 1'b1;
//	FL_RY,

///////////////////////////////////////////
// LCD config
assign LCD_BLON = 0; // not supported
assign LCD_ON = 1'b1; // alwasy on

wire io_dir;
wire action;
assign io_dir = KEY[0] & action;

///////////////////////////////////////////
// GPIO
//assign GPIO[17:0] = (io_dir)?GPIO[35:18]:18'hz;
//assign GPIO[35:18] = (io_dir)?GPIO[17:0]:18'hz;

///////////////////////////////////////////
// HSMC
assign HSMC_D[1:0] = (io_dir)?HSMC_D[3:2]:2'hz;
assign HSMC_D[3:2] = (io_dir)?HSMC_D[1:0]:2'hz;

assign HSMC_TX_D_P = HSMC_RX_D_P;
//assign HSMC_TX_D_N = HSMC_RX_D_N;

//assign HSMC_CLKOUT_N1 = HSMC_CLKIN_N1;
//assign HSMC_CLKOUT_N2 = HSMC_CLKIN_N2;
assign HSMC_CLKOUT_P1 = HSMC_CLKIN_P1;
assign HSMC_CLKOUT_P2 = HSMC_CLKIN_P2;
assign HSMC_CLKOUT0 = HSMC_CLKIN0;

///////////////////////////////////////////
// TV
assign TD_RESET_N = TD_VS;
assign action = FL_RY & TD_HS & TD_CLK27 & (TD_DATA == 8'hff);

///////////////////////////////////////////
// ps2
assign PS2_CLK = PS2_DAT;
assign PS2_CLK2 = PS2_DAT2;

endmodule
