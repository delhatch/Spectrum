-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mzL+OFHMZBHx5tMO4qfod6DiPuTTH0axA4QWYMTC4hjwa6l5v5Nw9V01wuLC+e0nAzio8Isd6R0/
38BD9sEI9YS63UzodbPOfGQtZPViEyQKIDQzib86lfAzq0kK/noBbTBRF81yDJyl0/p08ujePYgI
Cw5KcIC/ZOLcc3xqJGOefmApUOh6YJoDEM02rypjwdSOmtFUmv1w2KEc/mLQFtLtwTFhL8+CfHaB
4GAnXICw+vpnzWa+IeYP/IVFC6ElemqOoElH6jdKZ7CH9tG3A+EkI9cNjrfFekeVAKU3W2xRqNku
5s+WZPaQmWAuSJRVigmUHCBELffMOCmT+Y51Jg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
4TxiaZaPdojF3rjIStVsasnCjEEkNoaQ9MYxqVT8x/uLPnYO7MQCQmjAz0Vi8XY2Lm7pVl3TaOlV
XgtBfxWrcoDXBx7lKHsOGhXGJpm8hfNExnZYQ/2BrUgfmBsYg9Zt3g7BivyCDtduu0NnvD7pv9Pz
FY1vBHZ5YkFjCiFIui/iLnej5pezpSPipVld6BXIMbRTPZ5bV1swISPmHAVoWwAWzve6WsslWXOG
cTfbN6SXbzxNE9DHMpgyjJY3GY07guD4bTVOlrOWy/WFgbDgzYaY+PpKM3n+tdaNP59WR1LPT/97
Wy201sds8lYw9oB9gSl2ekCf7bgoL53X+Cfd4TNiFoxIGUN1dfcsjYg7F5EQBoJibVS/FvMfiPL8
FelBQq6fNVPGfa/XNEcCB5huUD4T+CAxzzmgDbBYa3Ce1H0sWepFen0m9+cnFOofgdtwmDbymSyA
Vcrrme4f3YOfzq0aLdEbzQDThg5pgAXFDZZ/X1FelmiJO/EUykVu2GuraUjCDyG0toTcCHJ9Ssze
NJ69egmTWcSHhdD8ns75K+AM9qF6bR7dcyhcaU8UOug/XXt9aJPr57v/g84D3tNj5XheqNkvO4xN
Rzhmav0msaWZN5JVtQrRynCxiWDDQaoh/YfGCejIoZFSIlOuIIQqDmtM30BGM7Wb2bWK/EXgByWC
908J3cs6jrNbDTo5uxmTFQKwecsECSsg5vPe881bX9cafIe9O9qg/AkYxpyxSRh0fL+2B6EY7NiP
pH8Aj72e3oOzGnHxJ/sdtp8psQuNltWIYzAav+mGaOxQO3kWsIhfYf2wvqXedVrbeUghY7tXqCPb
1OG4nayzsgvW5BGmErVWdT4OulDJb5fer4YGzZa1tvggGcrkZuu8CUOPOkn06R5XFzoXyO/ekPwG
AErZ7vQula++Vd5EiSHqNxatxuWCQm6OoJILUkGUV0EMDAM4rNqmHRJVgklxfOx5MYy7/WQDoOND
074c7La5qk3ZN9uAV4Jbog3DVK/q8CKgAk0qaZdZnfbMtH3ZeTI/BKk1eKysI8fu5vBkHA3FeZAX
LgUe6Ep4vV7T+Vu9y9Hi4wIvZ+pv6j4YhHC5dmw41BE+8fTIGorwjiukvtQ1zSAGSOm6Ow0pe3AT
gsmGy8oiW5zRdPFUdw8u0lY767yZgY/udPzxK19iyJP0lhJ+WDVFWsgs7dncfmTQf1WvgOWdQ98n
oHnaw4JmiQISihX1oJgseJZOvw6M3E6aZMBWeq7UGJv7XcLAKLYfyMTmgG/v+NOqMjU0qoK5AnGN
GAVZB2cTg7juzc+lj6zJEkwvI4jhIPFcjY3kkH4Jvsz+tHwweIHTRDsp4jFUHiz99JnTTfODur33
HhrNtEk1kJE6fkjvsDsPePzFWEF2omnsxKjLi/YZ1kNnTwa0rhmFqrUyMFkk9qYRcLjXJuPq+yqe
SprgAqWpynTrfVfsgjP3bCZ1LeWB7xttQGJoWl+YbNHnhxugkomsboZwwvxcGzmQVZNPz8XzSEUx
GWtVO26g9cB27xdaXMJ98AWVo7DEOVknfjmQyAZI1o58D6Q0mgcBCT0rUrlaZgXfP4GX5ygDJQq4
wPnVQ4BU/haDe04CSh7WzBjBNiDkOKyjmO9QxHPIR5oA8LwNCVW7210xAGHKavg9L7RB2fcBxZEe
yiIiqeicpZVp9qTW91TKrbG/+LaKDiLrUzJiVGASxpPvjJpPGEHSybPVUwVtB+VQazpqc/ZFZdUV
y5gCJ3duFyAI9grSoJKgZvmt2NkjTeuEFCRfhGSBReOMWYvFheDYa7nDeasafm6YY5UA8MgTX/1t
1mWuDKbp8A7JTssof9KamMLnoP7FdTXzjJMC64uiEomuniyYeswOVBr5gx3g4L7DGRdgnfNvgTZS
A0qwBNRDj4Hf28PlBGIfFaFTiEeXFeXelusXaBubJkX7LwdOteR/GZ3crk0VNtgpm7bUwERTOJNf
1QKtj4+3DaNyVe/0v40McPTve69iJyBYhTI9J4tmNPeInVSRO1sF8t56uysidG0Xf+b2RUOTSQVL
zQtn6VSujtDxMU8bQb/r7FQpI4y+iLmYtDQovS2DGkf8boUdhmrELL9tExO/LGGGD+f4y/NVS1N7
mjKSlECY38vYDbh5fIO8jbD4PdsporIMi504Y/0057A6Vrd6mA5rpb7hrFx6TAve+XgfA84pRtve
wWdBiowjyZaImasPeZHuTZxZ0LhKJHHrfv09gPuoKDQHCaRT6StMXmUgytTKVv0nttiFdTy6NLCW
0q1WjEfCdq+HbiLLZJoXhg9cjRxnYI4P13at4HRnDhbJUmlg/AlB6XD70+TxWVQSu4Yxj8vj3rUI
ngSuE0ibsCA5gMoOZF5O20vQQ+W5qKUtnkBXIC8H8VqkoPq9DXz4lmrEaBYd9xlqcrAnp6kIkIec
AjLLbc/++73Yj/z76ZyuXJvkvDTxjiSjnyl9SoW7DrIiJk005gQvJpzmx4uXcUacxnkMgQc0yJhy
/yzNHyrRN8L6KONxR/d2ndTP+kL/Bo/ix9lGeYIEXJFHD2xokKn8+c+qGovS+mPaGMg9KaBXZsFX
2zfSagFgPl6dPWB9P5SMxdkuzcYn2NGc+9dWgwGCrGdB8glWH7yUuueI/AepglDpjJtXqUwfgi0P
X0d1xk+ij8IQemPnW9NlMqz6xBaOUgvywuXLLDg88CT8z+Ox5tPTMVl7l47zDBhD6vrnZsZeTeaX
XKpRR/oyibcNN4dxFHlWM0UjgMev+B2qwZwGgJMIMxt7mPcCbG4hBgDyZr7CwxBqR+ZSDLm1yH2W
ROGHQJdUfac8JMnT7ex7FbLCMcReXn2xce4soQS8qRM10UpxiHap3qQtQwvgTxasCj+JW6pEuI36
VvdHRe7WMEmz6UoftRKzEcugnuNf3v0URryWZqxT7f3EF3j1w5k/mu971pt11uyGABFwcFSuTN+3
eGS0EKbYuZCSFu5K57reNtjQgiftbJ/ROoLgBPYdvA/0RpZmvBQ5eKU0ial0BipCOYPNHiWLmQbn
f4d+66V5hVJJKo0oP2OIon8c2BPpGfcw8MBrBqjBA3+G/T4AdjWsd6u1Xz4+HzJzndLPyG7z+hkb
A34O15dqkDqdBhiBGmfFtd6ZPztq+QphCtx1ofo3AzsnVMe09oNPIjyDlO9JcV1Jr42M7UmArLGv
96XSR3NNGVQ/QlOuTNsKXtpJUDEwGKE4bwC9PoHhiD0N9krkd2uRbtmbCwgsZgW1M2haGQrEozhk
Ni8SZgwyw1mUi2FTvZNvmdO6Kr7MVxAor5XkRzXCVYFKbgpaCx9cKdx64qQ+bF0BWwM+9T5w/Oa0
PP8gnuiWx9nkjOwC7cGn29fcHdmV4ggN+j67syrwXBIITVSm66TDjOxZWdM5jyIKlheNvPGSw3E4
tWzd68SnMI40JVUIuZ4+bDsqDraZ+E5tGXbWpWrTLYil+Xdy3RbeZg3RfoGThYLzieDzIYfFuzEW
+eTaoVG8D6DJYP27xmSBjCEDwJrbVgzQw3myf/Gyox9StSCtGVj4gq7vh+3GT3+Q+d3a/wwjNp8V
yB2Ue2mweSheOOh9BfBmfPqIoRcOAWBBKZlsrLErZTZCHjEaSE+cegYCdfgp28wlccOYhXX7HJ13
NvH8DsTLlpG4Vwi3y5eUaeVaSQz93fakb9kj6QpsobTwMtjn7bxnbDYTU5l4SmZV8YylyWDjiZIf
/xBlqMmEph75QZygnGW3JOx5koMh96I4r1zbl9WWXulglzloUIHUbvxmqFivxwuncoApOC3sVunx
LeNhULEu8r7ufXavIRy+Ywcdy0CVQ9qMLZug6/4xvQy0E+ljfbhPXmNJLc5zhZqPEoChy612gydH
vB1gzrN3uRIiXK/tiMwoFfyQulUHla/5PoxK+I9LRU5CUmzUp8OyQJW3gE+VsTC/qcDy7V4tSD7Z
C16Re7wpaAVe0KbkIH6lDiYz7u2XbEn3QHfafLMQ9ypDP8UovcxeQOP/KcxvHr1P5r/tshXVMU8U
fEXbIgGUfCXWrBTANYnOat6vXtCz0CWbDMuWglJkxmlhbNp0fpwI7l6NyDqL+VJZBHJbxuNfL+Am
5yj8qEGyzRExjfoyss/b4S83mPWx28UU5vJ4pYdx4pjvrtQvm2x2q4sATB9ftqN4qeYOFBojYuCe
eSkz7CuUYhDfBzSvvg522NXCm/v9Vys50GunLZmZBJW9EZq7t/xJkYGlvMMuebxtc0FjQmn11Cds
H452lmXl7sFZJtKBf5PiJ+1x9okepjkLPovPOWLpQBxy6xU7axAC7v6e1RmmPaGm1kyVe+futDMG
VhcIt+SehJB/FdD+O6XuP1IPk3qoz6Eq/z8752Trgnm/d1RNmz90iTMxVXXF62yi1YumM1LG5Xww
NCcHs/eW9uL2rrv3qzHvhBb+7ampGUI9BT2oCFlxuz+TkREczUv11TM/hcxMem6jWJov+72bNE+N
m1qzPMOvpJoXr4dqsPVTfTklTvutSTsbasCmwgwfYk+kQ3lKFdtPQNo1NqURVMJS7fl415pwvjct
ELGzhIuyOQWafH2jDItm6DxYqIugJkHjRxAggmij8PJkRzKeZJYSbi4bgfIC3sPtDXI+XJcsHY5S
h209hdApGg+5U6GoPYngAIMce2kIlbRrVJZqS9KweIv6BOafurMq/Y8P0NmrqgjKw2h5F16cqSRJ
Q3w7CwuswDZ0Av8m+qjwROwlajOa0NFuZERfFzkOpmhiH/lwPHnSCT+/xe9JP2GI7r5E9vdSt8vt
DCdcb+0qAmgKXbQrCLlBxuy3643qj91Jd12aJlRGgB3vzItZW/Uqe47mrwU5hBciE0XSNC8Ywp5a
0acKQYRJV59eqSHD0NX41LntsieEwPH4Kq97WeoAEUQ1YnScDJ+bljuazcdWbrqUH88Oo+s2d3JH
qmgujt5wED0AvCMm9Nmu9wGWeratiJ5a3i1X45kUob2o7LtFH6Vrf6nyXWzoatfdYbNVVZ4QF6OI
/NuUWgjQAZ2WQpQVDI33RXu/WeHw4QVOQz1fNNPTyEXuefiMV4loYBXKtvAtaT3rVkJh7s5MlCpr
4yNbPZwA1ZlllSLx6Dgc5eBYsS5MASbW3Jo2YvmnuI7okgZsJfSYqtPPYvTd+EWIV+jFTjzq13LU
W9GAqqx4gKOCZHS5Z2YZ9ntKCStyMZEMTDHH+4/Rzv+qoCSXNIIgtV5yYRlqpY7Xq887lf7+aONl
ZbqvteHNdo6kalLVVZVndCgY//f76UUhrIk57jUpA+/gIzvTBzQeqjpd0aZMtTLTl6Xhel65yeoE
e9YR+CeFaAQtHYZ/v/q0clb86kNrWmYs0iaxNqWCgeCTMIVJTsjRNxuZuG66x6eyy0IQqPpdkugr
P4IF8yBhPYrUYtORmeXDlvOfw75Tfh+fNeLHkulNw/10JZubFBJ/v5WwN5mYkPjyjTcKWQQ2LQNJ
7SNvIZgp+U1O2sqILpGSvv3PO94NFiX3VQeU3VPXMtEHo6NjQn2CL7EXDHQ9S/cYKhtTMALjDZJY
h/zn30U4vd0cL0KNoycMD7RPBZDD/8sAY5TG0JbfctTzx1yj24NGg3G9hpJJJFnfHq+cv+j9zxm8
jUfvg408/bun9In4SwxAKfWc2bAUTh39zz32e9XOCd+aza3uoFPhrxHWZkYj0Jk2u74CuuK2DTGC
t8BEW5bM6RzT6lcLHFexpRaWyxJRQvC4mFQp/bcjBzc9ayniHTbWHKDs8F0w0w9Qcxq4baIwBMi6
TjXIk+5SC83qkhqTjafdt1x8SHWrYO46iXpfQUp3vxtYNUHFlPixMn2mL4yatcEEu/hbVBhcUXzS
mvWoPJA/fV9Ovn4YAnF3+QQ52rz91Lmn2iAJgk3dFhtFPkr13Rbg2mvcDpZ7hsIBlwwgpYOWwJXP
V5mIGzJPhXCWhPiNSmMk1FTLzXvb50WdA/33B0j6EbbjSey8MOd10fykmjBpshcCQZWXx7BNQfPX
LCs1s6dxHK00Hl3t/V2EPOH0hB0yNB0fVFKK8UOYWmY8ouchLpzOStzlVOGJiobxCNk+++EDxbka
H1ADLeucFvf6KvXW+J9yypJfH/XCFYpdkg1WnN0bTFdvadsMqS4YlkNL6ewMh8jOEXsKmPem3e3D
hkdHMkAk01aYl1W1h2ziU3/tW16rbe31hjFOQbcLMIjiYd0yeVPKYKWcOnghaACpqoE+11z61amg
F+k50hPUmdCIDCNGvn3jvKxG2LfKKC2pFBhpRIgBAqlhiogJC9zs7k9eQxYmaYbV61JqKd9ctlJO
LA1v7F/2FfG1Hc4gQ7fiNYSNA4M16HrYWe8H+09KZ91vERz6/Z6Up2jvi9adUP6LV5S0uzGI6aY6
42DoCl26jPBqG0ZdLRMqUSNzKBW6ca4V/pIX9UgNnbfOvM+x9pArd9Srlow8TBMpAJAoHpKrtgVN
8J8fb/NcjzKq1goPflfufrsrntzQWD6YvTZfTw9r74XXmy0d6t7zqnnmN3cghSjsy4yiX9O+VVs/
YEIngxIhVZuxTKEVpbS2kJCZDkuCFEIcUJmOEkjryup5msNyEmN+PB7ZoPU/NZGrIhZxxAxcZIMN
4RL/HBYf/wBU052L4/Nn1ZhOJ4c368XF8kzftmR33Q/ViUZ0OMDuN0DeMSjq5v0HdAf2xeLNKFf+
voU327yxfOR75v0b68m5JxnQluPFqjUwPdWnI4C9JZSCcITubxreBAIoYBdN+E5aG6K0K+iuYcqI
Ov78K5vKf56n4nFGPld1NG+mZir/TOpuf+laK1lE3J7tMQ7j6eLcj4euvL4AAjEJnoq/EN/R+vvy
uFfv5gzEqkfT2+Sj64CfMQo6yYkloDrhhJKkdF776CizPA8b1wMbH95yTMF1PRW+Y/8aubxLllWt
ZvIbVJBpeTusOTpCs11A/rKxcIyBti5ijUJqgfiP3YEyV5O5GAPQPx/J4jP35+aNKfwRCsJSBpo/
zY/n/5Ke48dv4OQ6jFJXIkQkRo+qSTSMkzwx9m7kb8G1A2NBOjzaFKswfKcVoBGxA/EUQvsiecNm
p8euz/DzrfJQ0Y1d7DbKAnGBOEczpfobuR8r7sl9Nu3SaHifTiXFxaFLa8N86vM1luPzL9FE5VLm
3wQiu+WwZjQ1b1Srx7q9qWHGNO9CBr73pkazhU13HHao/eKyHCR16xmuE8bzYBAb9ohBl149P91M
zn0OhsXDYS9eLfry0VpGcfN9NYpNeSFxkbp7uspdWcts9mlcRpusCq89vjwsLjyW08Zi/ExR532R
tcnjFQOpZesjehS9zxaflBjRws13VZDWBC8sCMGg7ANceNzWXI4/E/ZoSOjvmgj1rRDk4YMN4SW+
DOnK46wHHHrXzdNIV1tvHjfO/68M8aF73tKTpoKy+a3QXgZEcwj6s1iL6bgX9JPCekFLbH59exGa
M8UE41SwWf1U2RpX4+IVYQL6yH9Q3FbHGaA5z8cyM6/+o5VZxLKipkJ8Eh7MeA8zlolhDA1NKDJa
aoiFG3iXgfk4LiXAXXvBRhL4fMu4IIc+oyMdlSCfACb9nogMaxGuO2HGKATKny3pygJjy31Cn3cd
hVHkkq1ZA8niwjTyh/jebAUVsWERmFaYIu3u4hmCJ28Ii1pscT3BprlMKMwmd1VyyvVJUbPcA598
BpS+jvFEPeM2vaxq9/lIWaBwc+D/TD2uHmwHPzEruhOF5IYFrssAk2YoOQbCqdgMAnAGXtsnp2gO
ewi6ZpdrRPYxvVSq9r1iHPuvYH88P2P67rZQA05OJTBIDrwSSVwm+nh4fYwnNmclF/1/qQMJ49C1
hK6paIU+tRQgXdwPU1+KuG5CoAAtLMbA8zRExKLxvwMdIjpPC16Z4YcjJ5rPQ+IkY+NEuwSL5n6o
saI7hyx69MEicPho+cAIMjMcyAWhYsOqs7raRdRMGmoppmwaiwR0RwCgbcT05Lb0rmPkHRN0V75h
9CjHesmYGUdgpi4RRuzM3u/i+RbZPKOfmX5W7b2ZEtx0i8auSeWrh/Vo2WBw0G6h34woaQ6YeFam
eAZJMhAUj6qsN8CzKlxC7ZKy66Mk9v3x6H5VTxGQX/Z7qJ0VJ2IIqBJc9fiIW8kEBehnyXcgOXYa
cST6T9mXG8QbtUgBHKk4VvJwTiGoJ6o9nmXZ6sNQhqBRv5vWNc4yweNcGeUFpsa3VTyCvqLNy7Vf
i84P/qpeR1WtUQOWZNxJNEptDRG6i2WJunwxJNudTQH8KXZQx9ELWzg1jXSlHWuoT5d6eBbDZviy
8UiaoOzAsqQFXwjU4yksz0xKx9ppOy9pskleak3rFjKBijoxPh5oYP0T398yHeqkEHX9GFybU93m
iL+Y3Ul/BxKqDtz3pjxKJi5U2qjzVREvLyB2/jJ+Qon5BkNPc/dz224kE1QTKBCR/8Luge3Pd8Zr
9v5fcVeiXQWNoU5vrkeSpF02BfkTuxuf8Ngn1h6e14SUPlpuAKv9Ffaa4a7Kvipwy95x4fQaBZ5c
Xz76jJnV5jUMH6W3WMgkqC3ANR1GfOsZ2J6jXdIW6YLiTAvetYirKK7NyNYRwh+m8V9WV2Xt3Fvj
30CKHXWeuw8WF6fytbj10wHEQ2h3e+XVMof6kmFvgiVZgAXb5+uIEFRZL5fhi0gcsK+GrJcZdWCP
p7XOTOEZL/FGPQqYNByvM/sk99YQsq5LfRrfhOnGxzix0PA0PKGAUnu1YAFRclyt6tj/HN3EgXJZ
PobNfqzZ5JV91JkN9pQZSi/eggzYVJxUQG8KryZlW3LOviSDbwzJBDCSEiBcsvF3HuYashLcIQPp
zCJkQIwg0v4csZzl/QUeG+kZHhN/8qhFsBdRYMOuhNWXcRoWVi2TWTwktEXmT1qfRBsTXd0YD6Sd
bJlM9X1qLBDhPwuO3MH1PoxBy5nBU4aJPG0DMoaaAQc318D6EmG7PG9780hXbuG51MxQDxR7wy44
/Fg/1hiD6JqbXmOKxWv/63DH9exKDhyiGin0mOI7dCCkWt5gGvHW9kXa/md3+4FVBIFd31b/n+ye
oM2dVWOPvFto+7cwL5oY1294NClqbpxh5K4le0rbB+N2IDvHHDfmHWsuR3KU24e0bfatS9rjXDhz
YbfLWeUSyG0atbORwCB9Kwe++RfBF49VIO5v0vJCR2JVDjXU823hYUB4ZP83jc7ITTTvdDomSm3u
F9j4nBP/vg1x1LNJGTvnIhtlM6PQWGH67RSP2M+VTL29AN+yKXww/uIbpCyl0zGfuFqbMQZIr404
V1wsvL7ikVvH3WJlci1Ks5xlz6ErM6DqGE8S23fCttZ7431Z37JuY7gXlr1WOIke1WJX9Rz6roNP
4Og7mbKNXFoQ8mOIsyr9HqKUQWuEsrtCUcl0qvf+yFw3loiAQDgjN4D7UFKVkKyyc1qBnpDInmdP
tsQCrMGmuIqKMPJkLJmrvFRtNEifbVFDGtuHlJCHXbB4MMbTzj1xvZVLPkFHsh0Dro8P5cC0mkyb
eJMg/QFlaxPFVd6HJZljMK47Zl6GHysh3vbn3Qcik08HCPjVBalz8YCak5B6ikXeb8qRDqyqvs36
uI9p6xdxvWWlPz0KFuHKTPNDKslujVu6nvMVrNeyMDdPIqL9qdjqoVBx2AREYJrFyxBtO0Ow2wNS
iXG3l1ZifW1mL3eFPCZ16Zd/W4G5s7UUqKCF0io1N6X6dMqUOXG2RZsquLOZSaJR5nbf3I8cRsmq
sScK8Czh0YeXJo1euWNcz0Pdvb7pHE25fKJfsDM2te9VGW5BnNFEEgnxJM5FRgcQuxKCqyR/Zg5l
Rev9fDianNPpgyI9WJoShuyP270h9+WbVhW/07urC7qoO4v1mG9MbVsPzJ49ej8oWrf6AvFZbVSv
Wp5xY/rkYb0hbHb5CQ1mUsU3wcHgH7hLrrP4k2XF+0SMeifSOaeCgFEkyz3DqhyVTbz2iy55FZ5M
y5IpZFg5tEmjtMPknMXWN4q5PljULEG36YAUn+8SbgXAatVmfIoNQ6CoGog0Bsz3tKyOxg4oY0/4
xmHxWXiqjIKijihAgyNYfrD9F6w9mRymdaL9ZZ7AP4PeBUNN/gYCONAsVJT7tFaLS+HX9uDiGxdW
g6VOwlBngzyzD8wfKgX9TpSX2VHHzmGb2tjOiWeRB4jjN4ah11ilHdVfw/ePo5Q1Z81fmGlS2zjX
M11VpDeZz4TTiCUHsjJDwHaHB+hfe+XV6/6RB97bpL3i5rDsntRBgWWQpl+wDt7fyoXKHTOEsnv0
drB5o38Vu9FmaVueE8MBouYk7EFkdPBjbK51JZGC27j8E/7yUWmywZB58+D6pqFxrA6yMQpeChcM
uzOyD7yWttQ1BIjJuPnUORPPkiCedQ49rU8UqdAHyh9xM6tjNGUx4eKmRjhjWzd7Z5n4URoomVFH
6hay08yboszEAGQtCtNNCz27BnI4UBG2ZbgKEpOHWX5d3li6kLcE9ZtSEeZY7Pbet3Re0Qy6yLHz
TfjAB6XtYrpM6hT/ZjwhoUSo7OQHCzW527/ipC6TcuijccERUbirqmFrp9HjIdy8FByGYxaiIWWJ
6/DOiPDw9oqoDZUhvjG6LVVrhs87THdMdBwoUbfIVT/f4Y7Mpcy5Zzzt8XtXv0q6kd6t2AzDAaXF
UPW3UDFzKmMF8HObxdZdBnDmTkiZaZ148tQU2+3GKbxkB+B7uNBxnTrIzRLnew44zBiXXWuiQI2F
j1JDJTJot/43ZQDBwFtylnsnyuxW6H3sdm0ToRLnYK+3Eh62EMk4PlIsPgF5x0WLaCMCKmtIUgZX
hNbbfGwYtjb1fNIbTssTG1IxqhvzY634SCf1y7t4E7Fx3j8g0YXGNXqfiYZri+IeZJO0uTHnJpPo
F/jQHbxHjejJ/kUBDK9x3Iv6Xg6BKVcF0UblvGMmjGcSdseFrKZg/uPRfRZutoav5kQoPpA+w0ZV
`protect end_protected
