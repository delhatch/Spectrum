// DE2_115_SOPC.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		input  wire        audio_global_signals_export_adcdata,  //      audio_global_signals.export_adcdata
		input  wire        audio_global_signals_export_adclrc,   //                          .export_adclrc
		input  wire        audio_global_signals_export_bclk,     //                          .export_bclk
		input  wire        audio_global_signals_export_fft_clk,  //                          .export_fft_clk
		output wire [9:0]  audio_global_signals_export_debug,    //                          .export_debug
		output wire        altpll_sys,                           //                c0_out_clk.clk
		output wire        altpll_io,                            //                c2_out_clk.clk
		input  wire        clk_50,                               //             clk_50_clk_in.clk
		input  wire        reset_n,                              //       clk_50_clk_in_reset.reset_n
		output wire        LCD_RS_from_the_lcd,                  //              lcd_external.RS
		output wire        LCD_RW_from_the_lcd,                  //                          .RW
		inout  wire [7:0]  LCD_data_to_and_from_the_lcd,         //                          .data
		output wire        LCD_E_from_the_lcd,                   //                          .E
		output wire        altpll_sdram,                         //                    pll_c1.clk
		output wire        altpll_25,                            //                    pll_c3.clk
		output wire        locked_from_the_pll,                  //        pll_locked_conduit.export
		output wire [12:0] zs_addr_from_the_sdram,               //                sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                 //                          .ba
		output wire        zs_cas_n_from_the_sdram,              //                          .cas_n
		output wire        zs_cke_from_the_sdram,                //                          .cke
		output wire        zs_cs_n_from_the_sdram,               //                          .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram,          //                          .dq
		output wire [3:0]  zs_dqm_from_the_sdram,                //                          .dqm
		output wire        zs_ras_n_from_the_sdram,              //                          .ras_n
		output wire        zs_we_n_from_the_sdram,               //                          .we_n
		inout  wire [15:0] SRAM_DQ_to_and_from_the_sram,         //          sram_conduit_end.DQ
		output wire [19:0] SRAM_ADDR_from_the_sram,              //                          .ADDR
		output wire        SRAM_UB_n_from_the_sram,              //                          .UB_n
		output wire        SRAM_LB_n_from_the_sram,              //                          .LB_n
		output wire        SRAM_WE_n_from_the_sram,              //                          .WE_n
		output wire        SRAM_CE_n_from_the_sram,              //                          .CE_n
		output wire        SRAM_OE_n_from_the_sram,              //                          .OE_n
		output wire [9:0]  avs_s1_export_VGA_R_from_the_vpg,     // vpg_global_signals_export.VGA_R
		output wire [9:0]  avs_s1_export_VGA_G_from_the_vpg,     //                          .VGA_G
		output wire [9:0]  avs_s1_export_VGA_B_from_the_vpg,     //                          .VGA_B
		output wire        avs_s1_export_VGA_HS_from_the_vpg,    //                          .VGA_HS
		output wire        avs_s1_export_VGA_VS_from_the_vpg,    //                          .VGA_VS
		output wire        avs_s1_export_VGA_SYNC_from_the_vpg,  //                          .VGA_SYNC
		output wire        avs_s1_export_VGA_BLANK_from_the_vpg, //                          .VGA_BLANK
		output wire        avs_s1_export_VGA_CLK_from_the_vpg,   //                          .VGA_CLK
		input  wire        avs_s1_export_iCLK_25_to_the_vpg      //                          .iCLK_25
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_sram_avalon_slave_chipselect;            // mm_interconnect_0:sram_avalon_slave_chipselect -> sram:s_chipselect_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_readdata;              // sram:s_readdata -> mm_interconnect_0:sram_avalon_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_slave_address;               // mm_interconnect_0:sram_avalon_slave_address -> sram:s_address
	wire         mm_interconnect_0_sram_avalon_slave_read;                  // mm_interconnect_0:sram_avalon_slave_read -> sram:s_read_n
	wire   [1:0] mm_interconnect_0_sram_avalon_slave_byteenable;            // mm_interconnect_0:sram_avalon_slave_byteenable -> sram:s_byteenable_n
	wire         mm_interconnect_0_sram_avalon_slave_write;                 // mm_interconnect_0:sram_avalon_slave_write -> sram:s_write_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_writedata;             // mm_interconnect_0:sram_avalon_slave_writedata -> sram:s_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                  // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                   // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                      // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                     // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                 // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;           // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;        // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;        // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire  [21:0] mm_interconnect_0_clock_crossing_io_s0_address;            // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;               // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;         // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;      // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;              // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;          // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;         // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_stamp_s1_chipselect;               // mm_interconnect_0:timer_stamp_s1_chipselect -> timer_stamp:chipselect
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_readdata;                 // timer_stamp:readdata -> mm_interconnect_0:timer_stamp_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_stamp_s1_address;                  // mm_interconnect_0:timer_stamp_s1_address -> timer_stamp:address
	wire         mm_interconnect_0_timer_stamp_s1_write;                    // mm_interconnect_0:timer_stamp_s1_write -> timer_stamp:write_n
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_writedata;                // mm_interconnect_0:timer_stamp_s1_writedata -> timer_stamp:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         clock_crossing_io_m0_waitrequest;                          // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                             // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                          // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire  [21:0] clock_crossing_io_m0_address;                              // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                 // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                           // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                        // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                            // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                           // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;             // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;              // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;               // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_read;                  // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;         // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_1_lcd_control_slave_write;                 // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;             // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire         mm_interconnect_1_vpg_s1_chipselect;                       // mm_interconnect_1:vpg_s1_chipselect -> vpg:avs_s1_chipselect_iCS
	wire  [15:0] mm_interconnect_1_vpg_s1_readdata;                         // vpg:avs_s1_readdata_oDATA -> mm_interconnect_1:vpg_s1_readdata
	wire  [18:0] mm_interconnect_1_vpg_s1_address;                          // mm_interconnect_1:vpg_s1_address -> vpg:avs_s1_address_iADDR
	wire         mm_interconnect_1_vpg_s1_read;                             // mm_interconnect_1:vpg_s1_read -> vpg:avs_s1_read_iRD
	wire         mm_interconnect_1_vpg_s1_write;                            // mm_interconnect_1:vpg_s1_write -> vpg:avs_s1_write_iWR
	wire  [15:0] mm_interconnect_1_vpg_s1_writedata;                        // mm_interconnect_1:vpg_s1_writedata -> vpg:avs_s1_writedata_iDATA
	wire         mm_interconnect_1_coproc_top_0_s1_chipselect;              // mm_interconnect_1:Coproc_Top_0_s1_chipselect -> Coproc_Top_0:avs_s1_chipselect_iCS
	wire  [31:0] mm_interconnect_1_coproc_top_0_s1_readdata;                // Coproc_Top_0:avs_s1_readdata_oDATA -> mm_interconnect_1:Coproc_Top_0_s1_readdata
	wire   [8:0] mm_interconnect_1_coproc_top_0_s1_address;                 // mm_interconnect_1:Coproc_Top_0_s1_address -> Coproc_Top_0:avs_s1_address_iADDR
	wire         mm_interconnect_1_coproc_top_0_s1_read;                    // mm_interconnect_1:Coproc_Top_0_s1_read -> Coproc_Top_0:avs_s1_read_iRD
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer_stamp:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // timer:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [Coproc_Top_0:rsi_reset_n, mm_interconnect_1:Coproc_Top_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [clock_crossing_io:m0_reset, irq_synchronizer:receiver_reset, lcd:reset_n, mm_interconnect_0:timer_reset_reset_bridge_in_reset_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, sysid:reset_n, timer:reset_n]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [clock_crossing_io:s0_reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:vpg_s1_clock_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sram:reset_n, timer_stamp:reset_n, vpg:avs_s1_reset_n_iRST_N]
	wire         rst_controller_002_reset_out_reset_req;                    // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	Coproc_Top coproc_top_0 (
		.avs_s1_readdata_oDATA (mm_interconnect_1_coproc_top_0_s1_readdata),   //        s1.readdata
		.avs_s1_address_iADDR  (mm_interconnect_1_coproc_top_0_s1_address),    //          .address
		.avs_s1_read_iRD       (mm_interconnect_1_coproc_top_0_s1_read),       //          .read
		.avs_s1_chipselect_iCS (mm_interconnect_1_coproc_top_0_s1_chipselect), //          .chipselect
		.rsi_reset_n           (~rst_controller_reset_out_reset),              //     reset.reset_n
		.csi_clk               (altpll_sys),                                   //     clock.clk
		.avs_s2_export_adcdata (audio_global_signals_export_adcdata),          // export_s2.export_adcdata
		.avs_s2_export_adclrc  (audio_global_signals_export_adclrc),           //          .export_adclrc
		.avs_s2_export_bclk    (audio_global_signals_export_bclk),             //          .export_bclk
		.avs_s2_export_fft_clk (audio_global_signals_export_fft_clk),          //          .export_fft_clk
		.avs_s2_export_debug   (audio_global_signals_export_debug)             //          .export_debug
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (22),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_io),                                            //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (altpll_sys),                                           //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                 (altpll_sys),                                        //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_sys),                                                //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	DE2_115_SOPC_lcd lcd (
		.reset_n       (~rst_controller_001_reset_out_reset),               //         reset.reset_n
		.clk           (altpll_io),                                         //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (LCD_RS_from_the_lcd),                               //      external.export
		.LCD_RW        (LCD_RW_from_the_lcd),                               //              .export
		.LCD_data      (LCD_data_to_and_from_the_lcd),                      //              .export
		.LCD_E         (LCD_E_from_the_lcd)                                 //              .export
	);

	DE2_115_SOPC_pll pll (
		.clk                (clk_50),                                    //       inclk_interface.clk
		.reset              (rst_controller_003_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_sys),                                //                    c0.clk
		.c1                 (altpll_sdram),                              //                    c1.clk
		.c2                 (altpll_io),                                 //                    c2.clk
		.c3                 (altpll_25),                                 //                    c3.clk
		.locked             (locked_from_the_pll),                       //        locked_conduit.export
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0),                                      //           (terminated)
		.phasedone          ()                                           //           (terminated)
	);

	DE2_115_SOPC_sdram sdram (
		.clk            (altpll_sys),                               //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (altpll_sys),                                      //       clock_reset.clk
		.reset_n        (~rst_controller_002_reset_out_reset),             // clock_reset_reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_sram_avalon_slave_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~mm_interconnect_0_sram_avalon_slave_write),      //                  .write_n
		.s_address      (mm_interconnect_0_sram_avalon_slave_address),     //                  .address
		.s_read_n       (~mm_interconnect_0_sram_avalon_slave_read),       //                  .read_n
		.s_writedata    (mm_interconnect_0_sram_avalon_slave_writedata),   //                  .writedata
		.s_readdata     (mm_interconnect_0_sram_avalon_slave_readdata),    //                  .readdata
		.s_byteenable_n (~mm_interconnect_0_sram_avalon_slave_byteenable), //                  .byteenable_n
		.SRAM_DQ        (SRAM_DQ_to_and_from_the_sram),                    //       conduit_end.export
		.SRAM_ADDR      (SRAM_ADDR_from_the_sram),                         //                  .export
		.SRAM_UB_n      (SRAM_UB_n_from_the_sram),                         //                  .export
		.SRAM_LB_n      (SRAM_LB_n_from_the_sram),                         //                  .export
		.SRAM_WE_n      (SRAM_WE_n_from_the_sram),                         //                  .export
		.SRAM_CE_n      (SRAM_CE_n_from_the_sram),                         //                  .export
		.SRAM_OE_n      (SRAM_OE_n_from_the_sram)                          //                  .export
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_io),                                      //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_timer timer (
		.clk        (altpll_io),                             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	DE2_115_SOPC_timer_stamp timer_stamp (
		.clk        (altpll_sys),                                  //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_stamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_stamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_stamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_stamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_stamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                     //   irq.irq
	);

	VGA_NIOS_CTRL #(
		.RAM_SIZE (307200)
	) vpg (
		.avs_s1_clk_iCLK         (altpll_sys),                           //              s1_clock.clk
		.avs_s1_reset_n_iRST_N   (~rst_controller_002_reset_out_reset),  //        s1_clock_reset.reset_n
		.avs_s1_export_VGA_R     (avs_s1_export_VGA_R_from_the_vpg),     // global_signals_export.export
		.avs_s1_export_VGA_G     (avs_s1_export_VGA_G_from_the_vpg),     //                      .export
		.avs_s1_export_VGA_B     (avs_s1_export_VGA_B_from_the_vpg),     //                      .export
		.avs_s1_export_VGA_HS    (avs_s1_export_VGA_HS_from_the_vpg),    //                      .export
		.avs_s1_export_VGA_VS    (avs_s1_export_VGA_VS_from_the_vpg),    //                      .export
		.avs_s1_export_VGA_SYNC  (avs_s1_export_VGA_SYNC_from_the_vpg),  //                      .export
		.avs_s1_export_VGA_BLANK (avs_s1_export_VGA_BLANK_from_the_vpg), //                      .export
		.avs_s1_export_VGA_CLK   (avs_s1_export_VGA_CLK_from_the_vpg),   //                      .export
		.avs_s1_export_iCLK_25   (avs_s1_export_iCLK_25_to_the_vpg),     //                      .export
		.avs_s1_writedata_iDATA  (mm_interconnect_1_vpg_s1_writedata),   //                    s1.writedata
		.avs_s1_readdata_oDATA   (mm_interconnect_1_vpg_s1_readdata),    //                      .readdata
		.avs_s1_address_iADDR    (mm_interconnect_1_vpg_s1_address),     //                      .address
		.avs_s1_write_iWR        (mm_interconnect_1_vpg_s1_write),       //                      .write
		.avs_s1_read_iRD         (mm_interconnect_1_vpg_s1_read),        //                      .read
		.avs_s1_chipselect_iCS   (mm_interconnect_1_vpg_s1_chipselect)   //                      .chipselect
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                        (clk_50),                                                    //                                      clk_50_clk.clk
		.pll_c0_clk                                            (altpll_sys),                                                //                                          pll_c0.clk
		.pll_c2_clk                                            (altpll_io),                                                 //                                          pll_c2.clk
		.cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                        //                 cpu_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                        // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                        //               timer_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                   //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                      //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                  //                                                .readdata
		.cpu_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                             //                                                .readdatavalid
		.cpu_data_master_write                                 (cpu_data_master_write),                                     //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                 //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                            //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                               //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                           //                                                .readdata
		.cpu_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                      //                                                .readdatavalid
		.clock_crossing_io_s0_address                          (mm_interconnect_0_clock_crossing_io_s0_address),            //                            clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                            (mm_interconnect_0_clock_crossing_io_s0_write),              //                                                .write
		.clock_crossing_io_s0_read                             (mm_interconnect_0_clock_crossing_io_s0_read),               //                                                .read
		.clock_crossing_io_s0_readdata                         (mm_interconnect_0_clock_crossing_io_s0_readdata),           //                                                .readdata
		.clock_crossing_io_s0_writedata                        (mm_interconnect_0_clock_crossing_io_s0_writedata),          //                                                .writedata
		.clock_crossing_io_s0_burstcount                       (mm_interconnect_0_clock_crossing_io_s0_burstcount),         //                                                .burstcount
		.clock_crossing_io_s0_byteenable                       (mm_interconnect_0_clock_crossing_io_s0_byteenable),         //                                                .byteenable
		.clock_crossing_io_s0_readdatavalid                    (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),      //                                                .readdatavalid
		.clock_crossing_io_s0_waitrequest                      (mm_interconnect_0_clock_crossing_io_s0_waitrequest),        //                                                .waitrequest
		.clock_crossing_io_s0_debugaccess                      (mm_interconnect_0_clock_crossing_io_s0_debugaccess),        //                                                .debugaccess
		.cpu_debug_mem_slave_address                           (mm_interconnect_0_cpu_debug_mem_slave_address),             //                             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                             (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                                .write
		.cpu_debug_mem_slave_read                              (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                                .read
		.cpu_debug_mem_slave_readdata                          (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                                .readdata
		.cpu_debug_mem_slave_writedata                         (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                                .writedata
		.cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                                .byteenable
		.cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                                .waitrequest
		.cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                   //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                     //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                      //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                  //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                 //                                                .writedata
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                        //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                          //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                           //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                       //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                      //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                     //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                    //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                     //                                                .chipselect
		.sram_avalon_slave_address                             (mm_interconnect_0_sram_avalon_slave_address),               //                               sram_avalon_slave.address
		.sram_avalon_slave_write                               (mm_interconnect_0_sram_avalon_slave_write),                 //                                                .write
		.sram_avalon_slave_read                                (mm_interconnect_0_sram_avalon_slave_read),                  //                                                .read
		.sram_avalon_slave_readdata                            (mm_interconnect_0_sram_avalon_slave_readdata),              //                                                .readdata
		.sram_avalon_slave_writedata                           (mm_interconnect_0_sram_avalon_slave_writedata),             //                                                .writedata
		.sram_avalon_slave_byteenable                          (mm_interconnect_0_sram_avalon_slave_byteenable),            //                                                .byteenable
		.sram_avalon_slave_chipselect                          (mm_interconnect_0_sram_avalon_slave_chipselect),            //                                                .chipselect
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                        //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                          //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                       //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                      //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                     //                                                .chipselect
		.timer_stamp_s1_address                                (mm_interconnect_0_timer_stamp_s1_address),                  //                                  timer_stamp_s1.address
		.timer_stamp_s1_write                                  (mm_interconnect_0_timer_stamp_s1_write),                    //                                                .write
		.timer_stamp_s1_readdata                               (mm_interconnect_0_timer_stamp_s1_readdata),                 //                                                .readdata
		.timer_stamp_s1_writedata                              (mm_interconnect_0_timer_stamp_s1_writedata),                //                                                .writedata
		.timer_stamp_s1_chipselect                             (mm_interconnect_0_timer_stamp_s1_chipselect)                //                                                .chipselect
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.pll_c0_clk                                             (altpll_sys),                                        //                                           pll_c0.clk
		.pll_c2_clk                                             (altpll_io),                                         //                                           pll_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.Coproc_Top_0_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                    //         Coproc_Top_0_reset_reset_bridge_in_reset.reset
		.vpg_s1_clock_reset_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                //         vpg_s1_clock_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                      //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                  //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                   //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                   //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                         //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                     //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                        //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                    //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                  //                                                 .debugaccess
		.Coproc_Top_0_s1_address                                (mm_interconnect_1_coproc_top_0_s1_address),         //                                  Coproc_Top_0_s1.address
		.Coproc_Top_0_s1_read                                   (mm_interconnect_1_coproc_top_0_s1_read),            //                                                 .read
		.Coproc_Top_0_s1_readdata                               (mm_interconnect_1_coproc_top_0_s1_readdata),        //                                                 .readdata
		.Coproc_Top_0_s1_chipselect                             (mm_interconnect_1_coproc_top_0_s1_chipselect),      //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),       //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),         //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),          //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),      //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),     //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer), //                                                 .begintransfer
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),     //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata),    //                                                 .readdata
		.vpg_s1_address                                         (mm_interconnect_1_vpg_s1_address),                  //                                           vpg_s1.address
		.vpg_s1_write                                           (mm_interconnect_1_vpg_s1_write),                    //                                                 .write
		.vpg_s1_read                                            (mm_interconnect_1_vpg_s1_read),                     //                                                 .read
		.vpg_s1_readdata                                        (mm_interconnect_1_vpg_s1_readdata),                 //                                                 .readdata
		.vpg_s1_writedata                                       (mm_interconnect_1_vpg_s1_writedata),                //                                                 .writedata
		.vpg_s1_chipselect                                      (mm_interconnect_1_vpg_s1_chipselect)                //                                                 .chipselect
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_sys),                         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                       // reset_in0.reset
		.clk            (altpll_sys),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_io),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (altpll_sys),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
