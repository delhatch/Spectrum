��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X���_B�v}���8Z|���-�;�E�U��aP�JDQ�N!�������V�X_8�/j��m���\�|Ƀ`���Q-�����h{	@')bkyݜ�.�Z������K����,��h��\]�f��ʷ%���u��K�3�"ؿ.�b�3Kr������Th��t@��|����������݂ѳ��p	8����Wz�����N�{r<��2g����5$iK,��S���29�li9��Z��Dyu>��NRR��uΌ�}��佒�K��mZ��`�L`�47�U���y�J�<�s<T��[H����Vn�C�'2�bR�
�\q����u#uO��F���q��ρ�_P��s�w��i7e�JSٵ{$�T�7�@d�&��1��Tn�n�:�h�g)%*�����Ff��BcJD�x�"��� �~�i��\���5�����8�~�E����V�ʔ�_�LSI�+LlI��sm����e:���i�*�%��^C|e�j/}"���êlI����t��L폶pRs�������
?l��b*x�~p��E5�܇��=�#D�U�FB^�)�j��N#�*�P���`(ߓgP�lw���Mo��W��ޥyttr!>��L�"�e ��d�'c.E*"�z�hX����?�Ƅ'5#cma�EN��R*�N,�j�X�K�	eJ��񕓔���%b@��������HԴ֓�ɯ���9{�C[i�CRf�I�hx�[*(8���:��8{�<�����C���6�jo�p�M��e�K_+�`�t�!Fc�9���$��0�~7ԩ�͏8/�`�ת��s���4v�;�sU�D�Z�Hʯ��X�E����v潣�xv���,ú�����Xx����T��(�۔��������t��"D.��W|��9�j�4�K�u,�m�����=Z��+c=�.��A-�n	��E��|2��h	x GU]Ll㷿��V�v"�d_��p��k�1{i3�~�|c���:WdS�|�R(��d\�[m��Pd)��$�m\30B��P`�I�Z�If�J�uo�?4e��Mv��f�7�;�[4�&V�B�Չ�)RR�����%��B��D@"b�xѺn���R��Ɵ�ˊ���7�2�0���&>xCD�S���b�s�����P�����㼥��԰6��f�Ip�!��:wwB��q"'���N<�y�v[����}Yl٬^����+����BNp4��H��%`��M���]�<-e!wϷ ��$�s��m"�:�}G+%��F4���?|E�akS��=��q��^�L�ɱ���<ɪ�q�edst��6�5�B4=y�T8�j����5�����&�P;'ɾ6�wi`��Hb]�4e�b��������t�w���j�BH�V!��� ��_����jKn�1�&�b��3=�R�r��k��"HI�J�P�לC@�G-9)��+�^�
֠	��~�eFr�6P�w��O�@.���Į�-���LfSX%Uؒ".�����Bs�i�jI3����`�J~{G����3����W��,��y��Ka�[: �GT������g��t�9�m���M�"�	�32��!�={y��,�|p�F�n��,V(x�=s��ǹVA2�������nt�~N�1e�xm���{/60z�$�[_�{�6z^���&�+������.�!�m ����6D��N����A`�Z�g#���=�*��WG�Ei+$x��1B��?����� Q7}��;�(�*���	��J�p0G���w����R>Wo.Io'o��;�m"(>
�oV��6�T07�:BB#��Ҝ�\'�Fl��L,������� s�ۨ<�{�/l���^�Y����<%���8�E,�g��vB����<�(�8��/��E�����^;W�%#��*F�J�Qp@u����6i�X�ݛv8|*4L�[3;�w6�QN�u����=�a�o���hZҒ�z�����wG����zf�c����ػ�~��3V/��[����3���!�\Cv��@ݵ@�Xǻ��G�@�'5���g� %N`�����>X@��>�!=����3׮�'U� ;�!���:��%.t��6��O�˳e�P�-ǟ�1�Ff .�O}"� _���a�,Eg�U7O��������'F�
a��L|�v[oU �<�um���G�
�np*��f���]�/J�!nRh���^e�VIP��2�gd+;K��}&�.!�Ԩ����B!'hT�da���}f�õ�.�R͏o:<H���̟��c�{M,�2���4�vs"�|��%�A�~-�`���!.��Ğ�ǖu�ڵ�h�r���n����t��E�d/��}�Į|%G���{G�-�)�=1,#)џ��D_����d}�20�������4�N��Yo�EJ�dYQ�������
["�G)L�$��ǂ��VR�p,]P+���+��G��CL����m���/���� �����,������@�Q���Aɠ(� ��R����M����E|{O������
��u&مֿ��t�ܟ�	�-?`�t�6~SF۫�����9��+i9�U0mS[��LԿ�%�J�D��� d�p�Q��>��w���H�� x�F�yʩv�K�`ܖ$Hg�E�BHE�;�iF��y�P=΄#�̝�ok�7kӥ�=����X�����s�bZܣ3}����,�/ad�tM���!IH��;c�A����`=���5'��
���5�4?���:5�aJ��������?���B2��%/\���'�'����n�	o�(�;H��4�6�m�p�͘�����Ux��)gX)Ѝ٩Q�l�g$���**�3��Ef��3������K�d`-Y d/&1�D�� JK���W�>�Q-�-7U�Ԕ���<��b}g�<L�쬡i�̹r��w\泴���6_<�~}��HPZ��l���1���ih�Ѕ�̪�A��U��a�=��MJ��-]V�P�#��G��t)bf���0���#��m�&*��*-5�̪���}���#�`� p<�䔥\̂��/9g���v��jCq�����=����O[~aI>��%�G�C��;TZ@��^ܚզ3�� J�Z+Ō�oY�76O\�H�5 �Vo3u"��~�M ��g)��U��̏�7�-�&�TVzΖ"2�FZ�sPF�V�#�I>y�p�W�=9|�g��Y�~�v�i��}_nxh�y0-/萼R��vpd���̳{j�)��1�G�ۂ�D�=�>����a1�ʯ��I9`Occ�^7�$Z���16	6�n^@��������>>M�Θ�'D�l%�.
��;^R
���x�������p���B�fI���=!�}(Ψ ����P����:<p$��I�B�Q����|PF�T����pb{�ʢ`��Sv��k��졤�w�ތw
ӊ��T�"�]�<�_��:EcQ�q_zc2��&ӹ�֨="ơ�,okm'�9M$'Gkȳ�KTr<i).?���{��p��^��*�ٰC�?���	t���.D���D�|w9�� j�H��'�7��fxH����;�r��9|C��dZ/Wk\@}����D��n����������*�(�v�Wb�?�0$}L<�j�'n���V�T��#��%T#M������h�etv�sql�-���z(O�2%��zN�9+|����������&�0hhI����D#L)dG��Vً���ǝ޴U��t(v�`�v�"��q�p[7�E�k�g<_�x�:h���O��Ӟ۹H�)у�����X�ʦ�d/9]:�Ն?�����Uԙq���x;1Ci���F����>jN^a�F����M���Z����릍���2���P�Fl^��<�@�D.0f2=�&ma�S^̽���\g VǊ�VWPuc+�B��
_��F뉩�va��=�7ߣ:��}C��Y�S��し��'��9E1[�߄$,U��5؏��`��H���U�K_MG�	$);s�Áxj�k�E���+����U�r���\8k��~/1�!�W�e�\*y���cǍ|�YD��ɽ�ڨ$+^{;�Z=��O�n��YD"���o�N��Rw��3�0K�^οXJ�z��C�ZE9+�0����d�l�)d�5���cN�ClF%���M�9�_ƌo~3k"�u�Z��#3
�O�D����F�'1�c<6��ڊ >9�	��N��cY��M᳒�����q�����ÌD(��Jwe�&2d��T����쐼%
qS��{�J��,� ܲ��&N���1�,���)B�r�����-Q�b�Ԧ@4%ˇ2�<{[��僨-7p�O�Xv���#��VI���24��ՙh���S��&7c�gYm���%���~�%W*q)�(�w �NYFb��*ov�����!,�0��*-��N���J����ٻBH�:e�5�\m�3�5E~ ���!�D�E��A���u\�GU�Դ�s��<冢JjK):d���z\�\�x�Ɣ�2�x��}�%���i�����/ �+��"k,�%�g��+�;�k���G;�����3O�j��q�;�U`\!�n��B8XT��ٚ/�_��G�|�Iٷ$��! �G�q�O�.t��c4�Jo��~*?�/�OPӱ�D�ˆ��zS)���g-ƈ�Ә�����2"Xr�L>�i)�jp�t�1�|a�g X�[�Li�����P'���TR�7z3�1�K���!��J�N��On2"��u�- t����^��w&��Z��]R���^e �\A�+��۬7�ы�w�\mt�j�ҕ$��4���h���LǏ�J)VղC��Q'�M~���ɶ��A��+��G�BR�N��GU�O$e6ɠ�)~P�"Z�͒XN���JͥS$�dsu!�ؗ�㺅��~�٦����Tw�'�]�u-Ӑ�&���a�c�kV�5�{��y��v�%���H��|	��G`	a���g����a���"�"2�\�=���ܿD_}r��)e�'�WMz�+-Vpח����5�z��(�"qX�!Ll����J�"t�J��3�G^F�n�[�K>��z���o�M?�S�N�3P߀$@@�j~_����'�)7^�o٦4�JY�$��+i6���olu�[Da���^>ja�|
ţ���� V� ?��q�g��Qf<W�*WC�ĄP$�ѽ��E�ݾʄy�h��G�D����F��@��?���q����v����d)�>�Ѩ��G���e�^ߎK��4�;"� XO��8�&T�n�.j��h/hŬ��(��܌�2��T�[%n��/[�E���,~��Y��fj��%�o��A��ȭ�G�@�%JT�! �ƀ7��B�b,��x��J��������B���	�)mv�Gg�s�:���,~M:�P���_����Wp��p�b�E�}0�7�D3��;��ƫC�#��Ǐ	��S���~��4��0!0�K��FK�pɵJ����d�~���Β#J��?Q��ܦ����Z�fA{��	��.[�����T��>cp�$�|�����@
ln����c���Ү3�l�>��%O�Z	{)�������d�2��.R:����&����m�1�nl�|cC�J�y�47�u�	>Dog��ͦ���?�,��3|�˸����]��'��3`�?���J� R��܀'2��󲗷���24�v
����o}
���&¦�9ލ���j=>�D�w�Ń&��U=ṽ\a7���}�3Ldh���mO���>���N��Y�`d)��$z��.��D��	���
9����S��,~��æ�͢q������ .���|'���& ,,Z�2��F�S��j�*�sX��F������ƹ�ړ��ٴH<�������i��u��'�սb�xT�_S��ӅG��������f�3r��3C�M`����Cp,���/���j�9|zF -G�-�%^�lָ���cN%�NB]r<!�V?4jJ�U����/��6fi�) K0 Ȋ����|��,%�w����EM�J�R|�^�j?0ze}�׽��p�G�������b����
J���^��[�og���G�'q=<
��z��.���I�.���+ߖ��Qm�MZ��պ0���V,Ҙ�^��ʳ|��Q�aZ��e6Y�����≟&�=����ur	�Ʒ��LP��V�����I��%�`8h�*NQ�+Et~g)�S%8�\iV��E�Ou�c@;���44��� ep]o��g��"o��|h�}�m!�zU�2,�=w#A�zdM�� ^�Vu-JWx�`�o/�%gQ�3�ߢ̅���2�1ko���̳Wڈ�g�46��M8G�J�}����]��i?����V9M���rܜ��0Q�p%�a�6�cڂ���>nAb��l���ܿ�u�Q�����1��;�V��y�@Bp|�7eX��ۀ"z�L��D�^��i��Iԗ��˦ZL�L�H�xS�eRC�
��	���~H�>��гa����)^�ˢ�^L?���A=�;��K��ȋ V+��}_k߭LQȁg�3?z ����@�tg��MSi�4�5��Լ�b4���Kz���Tӕ��-A4�J��"P�oh���d��y�u;�\tRU�*xQ���;�>��o4(GY�b��O��W� �o�d�[��X����7���S�)Pw=%J�C��	K�!��ԩ|S:2@��"a(���z2��h�!'����
6��a�1,a��y�����kP�S��3��»X�t�K�O璬1W�L������w�S����#�B�E��͌)�1�BK�8wh�xIv$���p������ ����誠��7�iP����5>���R�W��>�\Ud�9�?�0����"��T��|w��K����'<�6>ev��3E�&r�&����S�O�`�W:�Ҝ�A]�R�l�� ǫ������������xL��Ց�����|k�� J�4b�$�u�����U7TZ,��4��p@�t�G\�q�5�3@i�#:,�ݒ���=�N�7�e�x��-� �:<�c�4������E��C
�L��{A�!��ܓ8�Χ#7<�gW(�y��?yԍ�$��E��8X�`�;ZY5��n�8�o�u�K��Ӓ�D�����|����.w�E���������r��C��a�S'�ޓ���߱=$  lI*��"�;�Б�~F����k��/ۺ�����KK�NԬ�B qԆ����B�b	xSi0d���>$�{K��[9�*�]��`����ɥ~KH3H
+���lˑٟM� �=1�1�!(�W��J;�sy�x��h]Dlᰏ������T��;�S�ѼB��n%}s� ��q���/O���(��*�k3��
q�F���G�ڝ7B�a��Y���2�?qI�g���3�z6�}�g8�GL�W|{<Pu�M<��j5�Ŕ�:}�mMG����R>*�h$���X׊ݔ��KU_V͘p�l\¬Fj��[���-BcY����@��`�%�Es;-����
���y\�܇��L�c���ϩ�b5��g���+��H�K���^`C6	qd�p$<ˮ/���n���nl���O�4�T��ϕ�3�5q��6��9�0xU�s�Rw��ϵ"�
z����:���~��ζu�@=���ԠA�`�� �vA��Qm�|��a�Ù.�|M�Y)	���8��KI6�۹�vO��F��Zo�r����ĵgD*>����b��%w�-�wP���1D'!�E�y?��������� D������;�j�L�K��6�:z��LAK��j�	��z���&/�I�@�����N��%���E(.`Ԝ^�� �i5�xk��H��P[h�\x�/���̅Q����n��5��J'�z�f G�@9���a"��	z�l��|8_u��lJϨ�K</30�6E��ЄP$-�g�G�Bf�.Dh�q"ɻ�z;�8�E�|g�O�qk�إ
jA���r�\���;��Oː�QL�DQ��0,��*#k�8'��-�e�#�Ӗ)�x'��l��2�
38�Z3S��K'؝k�?�B���v�1���w��bG���#�N�O�
�'w?��qx	��e�'�OS���B
���k}��[�w�b�#����)�{Iw%Mq�/�?	aɂ�j�޷b���J�:֝t��Xϣ��z8D`bÙ�kx���)��{D=�J\r�~��E-U��	c������0i{���8%�|ts"��<�B�ӕ�b�2����Gn�T��CEޒH�[r�bФWҎ����W�v�P&�ںf��t�ԗ-a֠�B���sя���÷���(?;���-u�Įp�o^�!���R����F��Kr݋�����TN�oJ�\Q����K
��ˬ���Etѐ�%�ꏝ�N���a�b��?vJ*V�v=� �^7l�>���\�g���������i�@�9���)�p�E����y���<�%���ۣ�ǔY3]�hV�V�	�:0�b�� ����S�+��8;���E����5=���ʹ���~,��p�j��G��f���������W�%�����G��[�G4�p�����e��Ͱ&�v6��W����V�f�i'�"��u<��h� >�r���2�-:��r�L��t������s��n�t �����a�5T�����G�Fz8{�{xV�o����D5��˘� U(嶋z�i�����{M�:��4�.�����A�)G��!�P�[�x�K~b��Cm���i��-W*ܩ����O����4
���(�M=;L�z��+n�$�gF��I���[�8�_t�8��#����)�LWw����S��Er��Z�;�����je1�r�B�b�����"�0���*� 뇗�Bm�l(/�����_7PE�K���T-�� ) fK���`ڒ��Ȁzv2�1$#�j6=P�	z*�"��s�@��9�#��Dޚ+�Ї2{V��DtS���Ϭ���+;�٦0=+�2�{4��3�P��a����&-,�(�ۈ���W������뙰PB�����Y?�%�\��%x�\���9��Fp���a���:�����&F�~�u��`�k��;�����M5��R����_���>���*�Y!��K/9���!�ہ2_�3>�8��hז|��Ci-�3�/*\eV�ÿ0���ö���r}�T��ę�oo�ܠ�~��E�����-K&���F�|"��t~ꇉZQu�������!ƀ-�5�k}@���L��JOi}�){����h�@̗"JW�^fh�oW�a���q� ��z�=?��Tx��6J��ö`	:=^b�EC5��)o������Š4��j��Y�.�~kyI���Dx&�]3̾�h�q?r�E�w����T&F]әPn��7����k���{�D��+����q	��t�[d}�o]4'f��f�jㆀF�_�Y�#, ���3�`�=xӚV~��(�V,V���-��\��EEa��P��|o�1>�C�Q�$�7^k�o�Q[T�$���h��]���b|��4�� ��r*K��)�ŘF?�!�f�`v�;=V&Ġ�Z��[X�B_�4�ii�*c��+b4�OJ.�+�5�I���g�w�w`�L��p_�t��g���{����L'S�j�E�|�J���S�i�+��ۃ+r��%|>g%C"���-�4U}^��!d���XH����4�T��ު V�_��� +�̖&�D��y4����
�P&���h�Rq�9���P �����d�<��J�(qI]�&��o��^j�l��t%��O�(N���\����E�kO�����Ԙs@s��c�0��'x�]��x���E�a�
����C�wg�I�����2紪�a��zH�8�K0�>%Q�8?��#�q�:��D냍�b�l���y�����{l�k��ǁ���AF���U�*3���
�,�:ZX��\�"n'$�:[�.S�.ȥ��m&m7����n\f� oo�Z�y�1�N�e���:NѥBho�s@4����x�����Z�u��݃�"�s'�~#��S����_�Z9�V����w��vL���Zm��Ju����1(s~����ę0�,����S�Fv�3�l��@'��{�c],�l2��Y��O1�m�{w�0B��	3�֥�q�;{���j�VP��v�1��u4�G��w����'F�hۻ1d�B�k��vf,=%�I�3���d�G�����t�m�m���$��%?�	���W�7��`nVk�b�tk��"�8���rl��8��^}(,ƕe�$�E��dZ�����(�t�ρ�OK�0Z\�(��r�H�e�[����^ޅclG�Bx�!��g����8v������&̿���`k7��(�Y|Oò��&ث�� 7�%F��m/sC��U&�DA��q�
��E[�-�Gi��S#T��dK���dɷ����3O�|U��윇]��Lj�@���F�eb��6�X�UMJ�u� J��5OF��۴
,�y�ۗ�X��zy=�㙘	U�}��7���\�ޓ���B �/o���?���l��M�����%
=P/
Cn?:�S��rCj��oۿ��;b���iջz0���:��e#n�d�ܹWؘ�1߸h�+[C��nD r�I{JIY3�.��l���1�f����>�Q��	5�0�<l��}ĸG��)�Q"��	.,�Zh�|?�S�e)W�c����b�s>��˫4cX�3����)V��䭞�xNx^B��NlV�G�=�H�����HCû�͠ꀋ*��5�P(xM�U���ɻ����R��P��Ʊ$IJ�2��J�V)Q?:���O�B�b��;1����4�:f.������~�m|����Yک^�*�����5�>�Y�!��^C��NQu�s�J�ӯ�{��O6���2�� kI��f����T{.F$hOs�b'�*�I���"(��v2JߎP�e%�� �ʠ��U��y��h�e���k�;RԌE�`Z ��"���$R�f�Z��I�qm����84&	��Y謵$k��ybP"D7w䜴�H�.�F�_!|��ڍ%uy��|����P6���& dT`E (�c�傽����qi�l���L��E#
\|�Vlγ]�8U%��Sw�/<*s�v����ב͓�T��}%��c&+��5D��=;_��;;�������(Jטm�ZB��~�9 T;�,nO@�[ϙ&+_��64f�t�^ɥ@Y/�/V/E���gP&��ĆL� �=��U�9���L��r�ɱp�b�x�*k_�X��I�"�����z�m����px�ﮨ�5T�o8��ꔴ�؛��8r�m��C65�3�ɭ�& ���>�����@`F��h����$������]�M�a��� ��+..
���� 4��Wmh�Z���ܳ$�/f{��b��]�n���1._�j�Ī5K����<�M#�B!����,%��{X$��w��ަ�-�'�4�~�����Y�b^~�~h
u/k����`a�q_��5i����v6����{�Ip��C���Ź�@�T92�Xa{p�ŏ�7�7�<���S��w�Qrf����� ]�rqi��qY֭%���{`_�Z��N|�3�uH>>�J\s���@S���k�ի�g���*K>��Wy3��0>f����*uqx|�}�-�z۬��{|d����kǽ�b�Ke�i��
���jy��!��x�,�����Z۲����h�	�C��?���+�R�ތ��e<��(6�Ʉ|2H�"i��Uw{/sT��l��h7�U�P*��Dg4?r�Woc�O���l죎βf�jGV"c�醙�n}�)SL�<w�C`�����H���~Mo��RTE�o):�P�NV�%~m��l��DD^���;�ͭ��O&>i1a1��o���X��:�YQ���F	��p�����S���Rز^6��_y1�}ӽ%3�Q�q���v�x9O]Z��?�ʅ��d�9J�&0S�t�PJT�a�Z�q��YB?�bA�%M S�3j�Sh��������f	��~����\���	P�n��&f�7�ɑ�gD<� ���3(�>�f�+�)	cR�RUi�.<��%�����˧
��t�A����g� �Dh�z���mY���|3#˿Ƣ����K��Q�	_1����3�a����g�eh�H����pdP�,t��ca3���T|_��^��
Ahxf�dNq�2d�-V3qy�a��P���ل�T��@a3�?ʸ8$��S��o�oj8m�G�0�q5���%Y^ F�!���l�g)�)K}q2T��� �{���֟�C5��rϳ
�4��*�)O��엋ZC�v_�T�� 8�o6�:�_%���?��?1�$,[W m�V7���B���ih��7�>"Z/�pG4�^
��][c(C-�b��4��Hyc"�p���2>�|�J��f��o���H�����\`��G�Y��1��_�MD�㐚!���)�k^�����♪�4�RFj�(�*a����W3��ݛ&��T��s��$!�߰���u���l�*�C7UZl{�Y(��_��.�l��-"�0��ۖ"��5��?#��3H^dl����Bi��0��0���	��О�=�o�N�ʴ+�̄	��)6�P���ŕ�e>ƿ���hz(���Σ�\�<�A�U�yE܏Fhzz��k�j }ê(������DD:ZB�{fm2v���6e�%�0�ͫ��A��q�,�Ŝ٫�& .�ܕC�I�b�x~ϖ���`�
��=���*��t=hI��j2�p1����N��5�FE�������h;ވ2��תJiBE<�GJbtBfpf���	��f�T�����ac���ȏD�5��ږ�t|6_�H`|�����70Yq�L\����B�4{�L`�u)J�ß�����%W��]�Q:0#��0fZ�=��T	{ �Ơ�$�<�����Tjߺ�l�����tƪ��@�(��,NH�M�L�%���a����V"�\����@֌<�Os���f�+p�+ђk��Pt�zL~��fX.�V2G�`tjPą����ĝ٘���9.&����չ�C��ʹ�xv!�*�X@����rk�~,���r�̯�	��q�Z��r,�2��%����"��\�0��N�1�Ɵ�lXVM���ZVغ �Q)������m��Wq�-�n��z{���C���$�}�89�B�d����Bm�6G�I<7��J[X���M�Ii�=�A�߅&�U��Z`��lE��cƱg+�Z�A�����h^2L6��`�M0Uk�"#�����<�J���Yg>�sl�^��-%�ɔ4��o����-�<��ژ�*���۽��nbD�d�{��0�@��ѥl�<�Q���Tk1��d��Lg��тr��:A�j�B̹���|�XC��if��pŖC��w��۱�
���η�,0�`Q3�����y����P�pC�)"�%����D��O�lON�z���I\ȯ_��˞nY	 �s3FU�-����C7�)���m�H�⚉k���2j�փJ�w�?���V�S�
��}�m�E@�ia�����/9�_	�2�[���ʃ����jou�}��ܮvϑ���\צ����*����_g�k��Fǜ�-��F`:��/o�uW���Q�h�ם1�1�p�Jc./�t?0�J5��Y�#�ڕ<�z�������B���RІ<��(M�T�.�����4�%tu��d��s�)�i�\�%u��\�=ɾu���k�O9���;5�����0�BA�H�G'�W�ÀO�w�)�
x����*Uq���lF`�u�䶂�����
{jf��[O�M�}�IqF����Լ���o��>u�>�F����b�5d{�"����|��C
c�E�X�!�J4S�2}!>qp�3%�2��_	�c4�C��#A�/U)�E��W�"q:�^�vI��B���=�Ѵ�f�W]]fH��DCv+bև�m������+��5�uɧ����{��)�S�n�������$���=��f��2��4NٌTj�v�-�lP
�^�Qv��WJ���U���D�I�����C�'-e��ls�>���᧹E�'��kL��zt�Gp��i�z#���*��*F��p	Qv}P)�h�_.i�]���E�-���n����p�
V�g�zw�@,pYtMe�r��e�B�g82��LE`ic\��z�պwKQ?8���W��.�L�Q�Wk�l�IAL�@�ᚱ?�1�>���,���j���&��P�6ă����Q��6��L��`dʭ(C�d�؛~E�8���I?9[2�݆�]9�U�y���]��tI���\���8Ɏ
o �|T�`sD��D�MS��Vz�U��T�y���nw�F���@�e�{��Xl9��?���U�-W�t�<�;R2쥠���J��i�8�-���F�'a�Վ��l�Do���3�Z���b�"������ɼ�B�\R�ܚ,�W���H�h0��m��i��:��N��=;�/�F=�����Д����@!�_\�]��r���f�p
�St�k�
z)Ba����rn�go��H�Do��Q^jb8||��G��&����r�D�d�&��3�<�ϰkL��r�Q�ݔnW�cu�(b�겏8��"d�%w-W1O��*�����xu�c�A��v�@c�Y%��K���Zm�Qࣨ��=X�w�1�{�!��]�}�#7<�Q�����)L�M+�TQ�N;�e>zO޺�?k�NCJ�����WUO���H����.)�T�+��u��.��,��ݲ��pM������E
�癧��0��՘�ii���,������ӽ8pT`�=�O2G�&J�j�M?�~ H������oG�0��h�;q]
y��&�v�x�i���V3c�#w~=\����
bgO<B��!͔���z,~E���P�S�4_ӻ��B�a�kT��������m���Z�Q��T2*�3��-�$7��T�@�u*��>�kY&k���9�H�����䗬_�S�e�f��'�5��;��+��'���-mF(��a���Jx2����8q�_�K����d�C�*e@h�A�#�ZK�Hyi@ma(kY�c���/h�\�ۑT�𪗚|�j5�pN�E�5��Bd*)����2B��0y�L1`��ў_�d�uCc�������1K_�5`���]��Ɗz4��4���*���xB�0S71�@��-8\���R9d�2�܈v�V�靍YE�����^|~��_P�˭��p�|�=v�پU�iE��R5��bs��\�kx��F۷���"�ǯ��ŝ�U�,bH�G��V��> *6{f㕄�����'��~�]~���'h����\}r�c�H�	�[w��1���r9���;^�S67�'ݐ��Ow��}�h������ju��qK�o����dk|��Ճ�ή���g�^D�6��	��$�K�I]���*d����U��ӣ:	6r8�T���s̈���g����'~�k�-��\J�g�u���HG������e��-�H|(��t1�=�$�2@�ԭ<��Ԍ��1z�1���O�}h�|Tտ�"��E2�sq� ��\�
|��y�����9��7��`{�(����׽8"���M;R�����,��J{�0�=o��$�<�ȱ3!α�gK=d�#��6p�S�w�G��u��������nDԢ�6�w&z�E��X�(DP4��pLN��:�RQl%zv��>w
ߨ�(�ݍw9>d��<5���Cc�צ��;I�L+�,��h}�P��.M���b��\�jn"�`��
�tH�Ea�V���9jp�/e��;���A��%7}���f�`���p���M��,�'���::�6ԋvO����b��Ξ��υ�Vv	�:�}ba	��u�^y��TSz��-g��(�1������� �ė�x�]����>d�%鶲�x5������n���<���iv�.��#Eد�~#Ƚ.� 1� ��ԯ, �����2l壤�8Uv�t�|���$�<�lc��x؋���:$�� ��4�"+��G`�����ݝ��vX�Kwm75C�}����Z�ٓ~< ������-İey?�����=_�ʃp��؍���ѝ���v��1�9awՔ3�!=8��5��o|���x�u�񒀠>-��w��Rj�Vڱ���z:i��9+&��7Bw=i'�=bS�SiI�㩎��y�֫`�6ZG����#&	3Kj����ă�%�gԚ.�r��h��\P�-���]��A���Z��Ha
����H�2�o���yT9���I&�:Ǝo�����:5����Eɭn�����`�D��P�KQw+�9��$���d0g���\m��H��	PA#���̓�ͨ�D8�b��;o�ɕ�A�;��p���, �i�|c�&��'OLB�N�п`�3��:9������ss	v�Ҟ�/&��N\G*^�� I.�C䢕Aj�VB�#�����;��wtiY�
�&��!�{)��л��j����=��F��Yl#�P�,�6,W۲ ��A�%#g|\��v����r�ۿ���O�������M��ǉ�-���t%"�r�������"�gv�-�k�Ж4�E���A���`s ge4'��K��'i� ������Ah���*�XA�(o���8��FևK?04��$�K����X�Y~���,wF	�/��rb��?�`mA6��t���>���M�R�K���`lmDUW�G�dK�z��,|�_�53d���Ы��k��z���G��tX��kU�ftg����;��խ�L=�[L����[�u~a�m�MUj����/����i�MM ����Yҝ�*TS���/пjO<d5�����H���XZz�h�r9��Oi��V��`���!�h�km7�=��[���=%�Ç�%��1���ݠ%��𝒛��4r�:O�5A�E���5�+��Zw*p LzSt�\/'_��_��LK�2\5�C��٘�ǡ|�	'�f5W0�)r|������)�II�E	r���#����~��G�U��z���7�I^��y���s���X�lW�T]�ʲ��#��n��@@	�(ù5�C�g��w� �vF2�N�"�@t��/���;<m Ѐ7V[��g��=>�e��~����2Q�b�}�:���2ԛ�h)}���^���:\8
��i�r�P����J�3֥L_�t��p���S̕�	.?F�k��'���=,��c�+Um/o������z�DNS��^l���t�6�T��� ����F��1�,� S*��EG92��8R���u�J�KN��Z�P��R1��Uh0����2i�`M�F��G��&�d�(�X�N��<�>=���eG���:&�"7$	��%��9���;(����<�^��z=��o�9(,�$+�s���ڽ͙�Wd�nY!�a�gZ�/EF���;{�,__�7`v���B��G�q��U�����t_�1�jSF+�o���ڦ�P�P�lm^�Ծ$�Xޅ�%�ץge���TP
Uy�4"I�#N�c"�Y��G�I"����@NĄJa����p[��Ŗt���X��"'��b����Xl��up�ԯs�X���^��2�]�M:����A��`���jQ�R5|�+M���M��%	�{��d��F�v���j�x�ǿ^���À������u�](3�\,e�G���M�>ϭ��r\ы;#�7�(O���@����*�]�$��I¬%h�	{���]e�0a1�,�S�4O�ԒK9����h!���6��AH�,��U�� 睊?������1a'���ؐw�7�Ttҁ�,%AŘQϚq�Gtc��k�����.r��͸�ƈ��˧7�N)��+ө�m�ۆ�e�;��qR�09҃����=N�/*����r���Ypu:<�7��B]���3l��O����
o�P�%�3Pw�˿�8c�L=�)�B�=)
Jo[f|�3GnE�g
O�����פ`��"}y��iO�]�m��Վ��6D�٘� 2S�>{<x�s!W�Hd!aR����OO���Q���P��2��-K�yfq+M6؟,wa2��V��]���۽��R��6��k&`."w%�y"w��Yɲ��֙��P�>6|����L�;N�;�W%���2��t.��})ĸn�n_Q�I6������R��.#Q�g�a��-A6X���	D�|7�~�d��ȴ7�Mѡ�L���}>�e]�L�4^�w�]���'��s@pPRgC�2����r��`�
#_�)!��I��=���x��'����&�ɦ�a:zy�3ϑ����%ф�\�q��B�,��؞�*��d�Q�<A���;��oN'R9=M�%*	����o�SUs�Nzp�.I������SH�)�
�I��S�������Mm�TV�;�i�3~

m�\��A�T�3Ě����D��X-�^}�c���Vwd���,���a�r�zu�fo��z������ʞsA�0�E
�?wpi]�+�r6<�4��荩�R�M���*8�$0�ɂ���%)�W��Js�po+�K#�l��Vl9b	Eg*��`�����F/���Q9/�F� ���������|E���{��x*V��qS��J��-�i.��B=�D��Oɵ~�T$0{甧,��RfK�4�e�g����٧��4�&:�a����])ɕ��<���ZlC729�~`ޞ�m]� �*���:x[$E��.������ ˠ�\���Lk-���m����<j�N=������/ӄP��|},��ֽ~��<��� 8�g�VG��v�J�/\�L"�$wb���0��n'|�JMѣK��˻$���D��`�S�����y����r�ˌ���;K�E�]�y<f�b>�"v��^֮��{ܬ?�MĊ�֨o�BT^+m�d��S�>����nAe��w��?^d�F[���#\~��b�^D�q$+���ٷg��׹�b/�g���2�%���6���=�a�bI���raΡ������(�z@����򢨒E	��zN�:�5�j�r^��.1�����+y(w(%����^ �Ma]�P�Ig�P����G��mɧ�1�ca&���
G0��Ǆ6�9�RG��eǪ��ZJ�5=A����ZO��1q�k��Tӻ�]j!<��'�^�}ޱ�F_� 8�֦WoD�|ݨ�	�$��<_�|,d��59d�jL~˥�;5��������N!��t�� ���r���|*��t[�S����8x��[���~[V3@.�"��}p��������D�C��ڔ����%6�pGb�.슲�e��YB�X�zV��� �|����[��ޘ�lOԛ1�'^hh�CmB���V���G?� ���k����Ř�J \�;�?�O�J`Y]l�q� ��'�QJ#_G|�9_�k��!���
�g�{��N�� |P�p���K�c䀣�.E�9!�@?��0*�X��r\�:�Im�f�zA�G"p�]��.6���)��M2U�H� ���n�eo�q\v����GVg�P�A�0n�nS��'x�D�?���<���@��W����RM���ت����vrʝ�	�{R�t�dŧ�S鏗���"w#��݃լ �0.L�6n��(���(-�L�"�-<{�Ƃ���y;��b�cZ�i�Q�Y<ہ;�%0)|<ZSjf���z����#��o�?!����~����I/�;�nRf9q��'�d�p6�i���hy����Zn���Y�|uYD�i�ӭb1Z��#QF8�B��[XV
�F��R&��x�}��k@+8�<3~`���¦�?����u �!>5���٨]�0`�W��]��zCm�o@���� a¿>�d���L9Z���wA�#6u�v��LXq��Κ�}��e�� ���xΦ��%=ITca ��d�g�V$4i���r�|X6��&6R\�Z�,�yo��﹫s9&��7��m���J�<�j���d�'��	n<�JR
7z���s�W�͙Aᛮ'&H��$Y���VU�%o�g�%C{e��ˎ#����ZB�9�uN� P��&*9,�moe�yM�&��s��a��h�aP�3_j8*�;���w"�ץ(�ҕ��y��w\�6$�.H9�GZY}�C3Fw���8-�'���ӟ��$(�6����b�rc����jU�`��,E��Ph�"����+Ћ�q̔N���-�YȤ6&Ȫ�Q����d�W�(8��z�=NS���N�in���eb�H�4��禐��F��&�=~Q1�;e�UÜ�6�Θ� {��ϻ�]If����-e��4ޚ!r� y� ���ڜo]7�M��Lut_!b�"��X"�a&N�/F'ib���%Zkl��{k����{nR=ag�(��&�C($�M8a��G��)���U�nt�~v)�Ȟ��C�,7��r��'��a�b�5�eR��;��j�~,�s}�$j���#�6�nU�T� �Y�o)0�*R���Z;���$CK3��
�@�B�����o�!�E��taI�� a9���D6e���ơy��yU������*��X������{�6�`�uR݆ofĴ�G��j�*c�T�t�>�4H��dg�V�Hd��/�w���>�J�k�"mG�f@u��Y��+�r�QԔ�6��~��B�|BᎾ��o����_Zl�i�Uδq��P+2��~*��ġ������� �v�M�߄Gj,��q8�%�:���B>��K*~�l'Q��=�V�r����E3a'��w�Y�)��$8<'�����z�Q�)��Ib+�u��E	�����Ӈ���n�o_]Ů-�Ir��jb0M޹g��{�?l��|�C��S��W��t�ah�a}�����^h����62�����?�y7��
<���HvO��j�ܓ߷���-�Jd�g$ZPb�_��;����~سO�� ?��a��di1�7��c台�%_{�����ˀ��9���G-"}M��݌h��侖�em�~�t�>rK8��o�����X�Fy W/0�޳
�T���_���0J���<d��Ȥ��|�&��,�&%&�k����|�C�+����gN�}:�&/�����~�����i:��=ʯ$�XC׀P���|+��Z�
�JU��(�F����id��~G�c�wim-`��m0���r�R�ώ�a�m+�Xz�麾���O)��\�I���щqWNL�0�'��(�7���?i)E 6��o�	V� a����ػ����V�e�Is"R��-l������\�|E[�f�><������Fbd��5��-ͳ;G��6���uz��ZJ/�T��"����Ĵn��Zfl9�\���k�kU��m�6F����|Z<�v�Q����;��U�[��zCha,O�ڷ��6ْ��k���Km
��n�O� H�f������@�:<Q��!�Ƕ�;�C.ډ��)�Y�l]P��(,���P �?ߍ{$ 76L-2�g�[�z^�c>��o��Hd���D���b��Oɐ�%��r�Űf���^ڎ1��ȹ�v�FJOim�P��Q�|;O�?�0��UZ��X0-/���C$R~L%j��pPf�
�>䪢�*�P}<w7]��ByxK��RR�s�ª��a��i1eF��fy��6
�@R�PO��v��r�:f��{g�"��9S@�{-�⠰��[����ԥ�^�9y�<��ä�T�k_!X�70���fo�0ı��Q+���i�&�����TrJ��`�\��o� ����G��P_�<�;�E[Nv�;�π ��إC�vO6�/@n�]�ﵐW�B�����t.��P��|�[.�ky�wAF������AJ�ӊ�p��k�E�r~�����t�m:ox^��eZ��n��\>*"�9g{�55��kpLg��x�V���d}��H|XR���]W�+�H?
���dw�� �PE�J��-��)��,�`��� �]�Q�bύ|-;L��ّ������]�-��Y߱�y������L��l!q\i3��j���S&��Q��@�K����]/�o�85��"/-r�k���o��K��+�����ȿ]UNZO�lb/n�����"@��bY��R����]GU>��{�Pu�R{[��uH4��_1����E�A'�R�/䱝wM�VMQ���g�F�wK���f︯��d��P}��+�t)��Ʃ_��`��V�I��kPkY��0��a!����5aO֔MOr����2I����=w\��}�p�j,*�vP��j���`�*�9���� ����G6y��a��PµZ�zW��o{�#P�����,���G1����.�p��K[)���z\��LJb`��-s�H6˰�>qm�p�g������~[rk~g'b��=�7���L��w?��M��nV}��`��m�?�N~7�=��i}�,�E���`������"�)^%�����)��\��I�"�8�)6Ajva��{�D��7�.���F�	_O����c|���&&���@.߀~��a�p'�� �s�!����:;_�q�s��:�0��Q�Mh�f�Ӣ ]g�>�,��4��׆()�⪛�Ȉ4���q[{�\�h�&��a�����0���v"�1���_}�#�Ð�����4��K� ���M.���(�xm5p�W#^}t���>�@�fa=��9���XR�_��܌ S0Rc>s�x�69!�#|)H%)w;#�ʇ��c�MM&�j���,�F�{w��l�2����7Zʯ=:],��
�o�P�a����$�PqY
Wr�p����;�d2Z�10$��Tm�����.��9T��!��M�i��h&�ej�zR�mG�5���W�4�E�dT�^z!�޲��%} y~�;ZC.k U]�u�7Fg2\0�a��܉����7�^�.�<���;%c�c���ÄԱ��d
@��mi���Iy�c;���l�[�n�i'��=*���c���k�s��:�,�ZW��{�d�$D�2]N6��E(/Vڵ��pl�YvY�{!�Z�Q(�)1��Ma�����MҬji����y���{:~N�Q�Q �8(�0��<�՗P)�i�Ͽ��W�y�I��.W�[��`��Ε^�D�B(֖q����c��
���o@n�Ďv��[C�s�@��N���ZZ�(��|�|�o�)����"�WE�@�k��p�U0�q�7_|�;���7\\��݊��!�R���I鶧�R�I����0����t˿� �k��$x(�.��.���4^\<Cf�����*Q�U��?A.��L���0�%�,:��7�#���xE�%?�����*`�]�o���d뀿'�CY��.�_�u�٫ͨ�;.6�h������5�x�-�m���IN��'���
�!�V��N���+�j��~�&�g?y)p11�ZL5��[�N!0I�~K@2�n�/z�7���(�V*�K�*�~����Y�������|��-��+G+ߏ�Su�����.{� ���%����F$��$0b�,��]��T�>~9WO�G�n��%�fE����ju�����E�'���#�p7Q׈ ��X�*��C�_2�i�v�`�X8zf�Ic�#�����u�A��m
!�#�4U�*�ضؽJ��\��lI�}����3��Lg9B��	�RyU�f@��g�V<�uK�adM?k�9.��$N]�t�(��<��t$u^B�A3B��/��=K�+�;7���9��/�H����A�Q�$0��	����<O"[�xđ�H!�65�*��p�v3�Z�ee��i�(<� �� A"���x��m��z���l�I��?_$�1|�(�������㘎1'7p�G�/J�x���=�r!��lH,i�B�V�Q|GB:%j�Oˡ/ �lӺG]�+*�j�'�p]��o�vp�0�;S�
�*��0"���Y2��x>":Q���mԎ9���:@�Ƕ���/���,tǳ��1P�M�1l\�P��s�b5@��6� �(/b����񱕘U$�<�^<=���T�2���Edl�]�`��\'^�
bAɅ���Z�����S�u�u���)�L.&�;��[m����YV2���S:-��Q�;Q�ǧ�8�H7��!/�(�`M�&��	�=��s
�����	BؚDF���F���$�Y�,�z�[��|�kVۢ=��^G)7f4�W7�n��A�l��r�w/E[©ѝ2��-(�H�u���q5{���nb�w���dF"�Ƅ������c�><�Hzi��GD���+D�Η�Po7��l4�Ŷ�9�K��. [s���E �A��	�k�%r�3�2�3��!��"��A��L��r�����D��*����:��}�tU�Wd�}�\�d*t�22F 	���Q{;1����2�sĐ�����[}���`�/�W�u�S?e�
P��n�9��X��vhi��v}�T����NܺqEr����3O�\����` 5E.��A��*JI�������c]N�a#�V��D]��d��m~���B'2W(�;k��-�ȼ���:P�=���]��Մ��A��jA=x��'0B������N���q���Z H??�%2�0�	���:�s��s����� �|����)��Հ3�;�k�8j΄�訊Ɍ��NR�:�V�q���
X97�{��[�Zf���s-�&J6d8�oǓ
&X��Z-���n^�^{��������Fgm
&mSJ<�"�(C�@?�W����-�5�����,� �������>����뽥���n^A2�L�i ��3���=��k�lG����!��x����\χ)��4I�|����Vo�&��~�x�7[�q|����(�t�B?���a?���L�7�7N�N.�%؎�xsu�ۺ��!����KT{%������|&�Ƃ�sW������$��u��|u)�3�Ea�X����W���5�ux٭��~��>�)����j(X6(��K�&[�A���
"�G��Z}m{N���
*4��}x�����@��,I&'x[
�$���0�(e�	�Ɍ���a �����o��P�r�1]wST�Sb��(�I����!#�JV�����B�'��G�� ��,H�(տ��1ĮR���� ;|�ÁTϓ�����0`h@9Ѯ�/�&Jm�ل��ʒ( x=����K�L
,�m��2>��g�pX��>jx��JV�P5��u��B�"ٶ��H�иZn�,_�3D��d�nC�X�',��1Tsq������@6H���b�h	�:��ŕrR�O��mwѿ~8g_+�w}��:a��{�t1���6ngݯ�L�փ!v
0�K�/�yAu�̄�=�r6"�b�=L�o"�.���`1rs�W��p��0�f+P
c�<H���zR���R��%���A	4m���d{F�E�=v�;���Aڤ���A����-U��h���b�:�����V���VB��#b�R�P�;�a�Fy~����e������@pƥLj���fiN���c[A�A]l%pR�\r��L�As+
���Y���/Y���P y'��X�{���\��ʩ�d�.O�������I��Tϫx� �����_ �VG��(/4֩}Hyx��#�)W�F$���.�Y<�)�O������O��1� �^-����w��я]D�F?:?9����[z���b�/],a��yn�f��A��J��2�������,0~g�Z��������S��v\� 6P	�Q�r��j��aQ���@��C�Oe����*:������|	;8Ǯ��m��Έ�l��B�=5��&A �d-G�pR*i_=�( ���j�r�dx>����oo|�]`��q�W`LH5;�ɒZ�����|����S���Gq��H��S	�#ۣ��Ը�&��:�$U�V9���Ó�G?qs�I`N��t߅��:?��u��S&ư����?�����$��_�D�j�F�`-IKWW�B芪��1/�,i_^x��p�AD��,�b/,l ��$t'����Kb���/���_���b�"֥n��~�O��w�����Ľ7�k����M�m��f\�J1�$p��N�A�#���`^=b� I#�z��q`0T�v����1�C����,��N4ٮ��g{�R�h5/�} q ��.����ķ��b>��+��mexD����D<$�˔���7���,�T����1��D.��,�C����_
��|4L![t�.�b*�j�f��M�YE�`��pj���