��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H������N݆��Ȗ�����}������XQ�ǔȀ�wu1eH��F �O���6���5ig�a%���5�Ќ6\�f����^ŶG\{���6��5	��p��S}��jO�@m]�;�ˬzgv��4�i"�d-Ψ�C��2�g�˰i����xW�2���g�~�E<�?Up��%����
���'඼h�{��3�ThE_pסsKVJ�`�jϙP��M��U�3�=C[J�D��Q���
#Ewe�ki<�R���͍\u�K�
d�i'z-m/�D�3
�_����h$X�E��O}/u���e�{J9�������	eG���#$����p:��)�Ί�Y�=eV�W�gmt�còr�Ó�̠]Zm zZ�q�,L�-�]95-���&9%[�կ�L=%�����QF*�?����M�3.���N��cؠ�=U��/�㾽�"b�o�[d��:��r�k
��5���3[(�}���)K?���C_����1���1��c�C@��K�;������3&묙�����E�gI/�-����}�6����(t���v7��:]8���w4�Q�R✅�S�E���_d����r��X����$��`��t�^��N�&�����<f�
(t�6A��-;fCv�w�q�Ժ�i�/��;��|�i�KfG6������
�Z�O����Q��	�6������A$��oϜ��
���|�A�s"���������+���V�W��,"�<��u�n�FkM� U�X��`V�+>����xc����VM��Ș�'����F��)����Zi�A���Gf1�DA!G�� @����[8����已'�\)\'^<��$h�1'+s3O7��$�Y�dY�)hk@����ɚ��V7�^�)���F�HD���5ӈ��k������ �w��xO]<C�F����.I�L��'(���e��`���Io������h1h�D�ú-Jo��3y���l�*$#ٜZt_#U�k��^A��H��,�ޚ��̽���]�4�O�8FC��b�ï' �zjw�`��c�h�ی���|�d�\ ���6�	��u�[�wⶀ1����<��yp=3�;(*�7g��9�����i�MZ��S%��ʊ�����I�v2fn�W��ĥ̲�2�?�����B�./E~v�:E�L��s��NY�ͤ���H=���"es�_1�Uà���+�{�Ci�I0T��V덫���Pm]���:g�����6-e��&֮���k��}�ʛ�/����2�`L�b�;���7�i�,H�
��ɢ�DQ���N�w�0yi����ӫ҅��b�hMc�e�d���5�fS
�������+�!{�z�TҸ9��^&�����K
���qCW���HZ]���hD�ʺ�6�v�v��~�M;O`i���rJl��_�3��C��s��~�ˌ�K�<,p�^��{��#|�rv�S���:�(�;�F��E+I;{+'�nI��"�K����?�,��>����ꞥ���Z��r�[&��>�L�hM��Z��l�:�E�	��
'�+5�j=��۳��(4u(��Nl�7І
�T�)A=z&����4�LG�7��<jUm�*���;�)��)��S`�eq*%������bSu5���5����t�u~�x�	\\տ2������J{��YOU2�%��Cu��d时�!�2���qy7Sy��i��8���p���ˌ�R��r}g[�	@Zi��kz5߹�=,���^-p���B\'�i�[��^J	+gT�����Y�G���Iz���K���o���~\�K	Ӓt���	��?�
���A���ɰ�ܦ-����w��[r�����Ǥf���j�ĢJ�#ٌ�^����r&GVCt���q���PFYz,�X�:X�2u�:H�n- X��ʹ�'�h���Y�s/��>{+��ߒr[C<>l&��	8�dLB �uG_z�-�:�b6��E�χх�Ý�y�)���#�Nj����|�/[^~He�E�ylRu(�G��X)�E��e(oxx�~�T�s�Gh�>�_�s�h
�*p�_�#����	���� ү�J�	��*D�*ؔ�� �9Ôr^A#S/6Cȣ�9h~W��rӘӠ��A!\V`���L�ţT ��y�6i'O"bG��Z 6���Y�����`��V�{�b}�K��>]�X_n�6���c���Mf_s^É6��f�)�����Қ����к,vh�n����49��K�$z�2�?l���(�����c�$��H�;I�ޒ�5N��CM�^RIf��ʭ��j؝�,Dh�юlҲ�B� vI7�]e�� 8\�:24b�B��7����@���<j}/ٵz��/ˋB��wg]@F�t2u#�&�/WǼ/yWۈM�6�R1��e?�A҂����,��P�<��@cͽ0f�����&��H��a�kb��Qq��9=?�� ��-5n3�=�':�!�&kF	�:8�X�;�c�
 �� _�N_8��N%�!e0��e,��.��PZI�AC�]�! �H��Dm���.��XI�.C@<����,�ۏ��؅�0.n�O�9^��\|����R'��[mG4�,wV���:ģ�G�-����w�JK�R�F���a�ₗ�J
�|�0�!�����Z߲��V��({����k8�%�V�Q���Z�B,� �Ӏ\8g����kh�tSe{[N������n滤|��2����h��'�5���+�e�6�vC�b���;�âs��y���s���������?#�5��~����'�e��������A�uZ���V�=iœ�r��Ct��v��l���fn\2��N�-y��c#���@�W
���~�M��<�Vx�M���k!���\�ǂy�����di}��Y��x�@�,s`W���b߆Z�H`�;Y]��[��0��U�ſ�ړSp|@Φ�X1R��.�d�U ��җ��r�~a$��[�t.
p9jZU�P�x�Sl{s�]�lc<@D�ĸ���`�j��8�s����#^�2ޔR�f�%��Nx(�<ޏ�.�Ҳ�Aꕕ�1,>�վ�V����([I�($U��h����9_nӃ�lѧS�\�N�4�\ߞ�%54,�j����e7�$�~�x6�����h'3U���+^�\����_w{�k�O�&T����V�'��$��q�цem�ۈ&V����ܭB�g��Q����H���X���{�Q�mU�U>�jB+_�z~�i]�j�o#���>p��~:�v�`1�g�6D#�������5#��G�&�K� Ov�U�LJՖ��fǿ�����^�F�LJ��0���ʗ��EF�6��|��m��� ��2n����ƭh\�u`��Ry��+�B���4��u���(~Bk�2���Ӝ�������t�U]Z��
T"��E��"�g�`�>5�ON#�ڇ�y�4���
B4d�sZ����\�o� ���
���Y�Vӕ���i��'�^�0+2 "T*/�Ӵ���`<2<)(��"�k[�:��	��?��<CW�_������9e
2���K�%b��x.S����������(�P�LeG*�T+�q"�g���.��̠����F*�"�T(�Q�x�����.�.[���7����ǲ����=*}���O�xw08�3�#Rg	��T�ۙ��e�+�;x����Gf���`��%SnL+~l���c��i�����3D1��B1��#���p�1��,ַ.�ヂ�ë�Ӭ��g�=�RH8�KÔ�x�
Kt�n��3�I�/�3����ԀO ~��
b�9�4�-I�[����	=�!�
r�j8���}Nݮ�
����+o�=�њ���q�Zh���7����X�E����C����a�݂�.����V	����<&h��������fMx��Tp�&N��p]���`��.��K(�=w�9� �;a���3?\�ǯY��˱��.K^�@���w��i�1����E�������_���1�d �ܕ�<] my�V�xP�<ݴ����F���ۇL�&Ez��<Í��8�--tm���3]ԭ�`{�K���T+��Oz�ru� �3�93���5��y&A6��T~��_p�C-3f.��s	��,0|�6���K�'}Dt�F
gϕØ�q�����A��o��mi��F\�V�3o̪�?�)AFo)����BD{ ��g�!Yg[�[}�7�Pή��ѥ�37y�)$�T�ؘVʦ��Mj�Q���ƽ�k�}F�ݶ����"�2�_I�@!-���%,VaD7}��I�Y���(�@d����]�@�X��ƬZ8�[�5Z+3���{�Fn�:o^vH�d�_��׏�Ld]����A������U#�u���yg����� �1�.�Bq(�W�2�J��\�B���X��j$+IÛBH��:�7�����fHW0���bN���;'6��@�N'��am�����;�n�ew{H�����0� ��ц9#!F�3��ө=}*sCF�2a7�ݣ�G/ �'��&Ȇ����4]���,C]h����z���e�]���tN-�����3t�d����P"*o��/ѫy�#��.L����l�jP��B+�<	�F$ݙ- �#GP�!'������9�� x�o	cЩ<�WYX�@'�^S!/�uTY$%��~�F3ه�w����;�h"^6����Z���rt������
�X�B��ѡ*��f��pX��!jۄ�!<M��O�����c�c�;�̋aР���B��FM��u�_�h�<p5��)QށE��]O��΂>/�|c���{D�*�:'��=�����9L7x�IW��S{'��΢�-r{�Y0E�����Ĳ;q�=|-�Z���aH"�M�g �R['UO]o\^��i���B�CN]���M�5@�ce5ã����F�v��f	n���N����	mPL4hO-ꄾ3��X�*��/iQ�؍&׹���ؕ�h�jz@�P,2����s�_,�DP܄�0g=�7z~�~�Dʷ+�/j� .0���r�=���O!��4s˵v��T����VM�^���	ZK�R��7~lC#ӭ�=�B�s�p�Gi��` ��kj�̤���;:�VA]ꍁ�b�%.+5q�����<.խL#j:za���s������Jm�^Do>�P��B"���+2R�9t5����܄� e����=���h����p��8=��B��������-�n���\��a\f� -���2�>AUC�ѝ��������g��-����I)�2%��34��̯9�05xE<v���Z�S��y��u$U�qi~�i�F��(;�R�Y���Ԣ%��e��7ڐ��V%��=�����2H�$���qPSx>+�<�uߞ*��]oո�����Y�k��P����>�d�`�o5li�5L4س����>"����@��F����o��N��Z�E�	L�\�!xK�*C��I9�fr*�<�6��d��f�2z8eA�aO�����N����#�P��JJ�%���ڃI�=�L��k[T�C ���_��=��,�Vy2�����)�@�pIU]tOH�p�x�©Vk�7؇N�_��x��䓳U��GX��̷����Q�*/�y�)���\��7_W��C,u�<_5��è�4\��C�M��t���{T��p(ɂ��+�V��Y_��Ɖ��\Ch�]O�,���&��<4u�h�`"��C�Ƭ��ly�QIt�D����嚅M�K"��Ȣ<}�G7B|g�G>���v���Zn�xa��d��,�![�Е0r�.��qXzx�E��g'ȡR�+�<�yGb�rF?2u���)'��eI|=:�i�H�f�w}��\���Lh�NPN߁0�(�mׂ��ڎ����Lh;3����|^���)NwP����o9�n�yG�!T�&C��<n�%�����㸉-~�	?@"�^ P��l�j\p�(�dE�4Dw�);��OM��_=U;wb�X���c="�X�������6e<T#"�|%�/�bW�1x���i�V���AB<m��a���c鲦�E�r��8T=sS:�i��1d��Aq3�C�7Zj1cn�M�Ǫ�݉_M��{\�,�e�i�+\��)ť�<�L��eX����m$�����u��7[��t�v��A�gv٬���g�����c$Pgʈ~��2U�6��-�Y����]�����G���p���׎��7����9f�-�����/K�8g�-&ي`9��*j�_#h��DF{���ߒ&����� M��!��i��^ �篯wfv}O�X�@mtw\�k�7��l��ls��
p
���[D�6����7j�w�0V�>�8��8�-f�CqVd���STk�g��I9
m� ��;o �����y���6|ض�?6N����`z��
ۜ;ǵ��V|�2 ��Ftߩ'���M-�z �(á<�0�E�L�N��I���K$g���s�p����8�o�s�����J��v�!�Asb�l;��ո�N^݉= �f_Z#�)N5&H��ߋYD^6H��Ɍ�TAĆ*<{BM�z$�Qu�4�������|��k�M�q�Cn��ѭ�-������M	��A�΄��ϼ�N��}dZwz͏�>�U�ǉ�����:若�%	e��ӹ"Vr�	�N볆��A�#����+�c�@�;�%��)�(XY���1�t���ɁJ���t�o�Y��0����\V�^�Ti:ʙR�j�S�ڣ=$��ub�wW�9Te�^�{�T�1n��U���k۾$em�tG�K^� Չ~rPV+�e��3B�ڇվp�|���C��m��7$)k�\�O�Y���|2�ҳ�5�p�,��X��]�C��}���ޖ����\�i@>?2�)�E`������z�M#������ɟ�����pimR��9,��]���Wa}V�3����!`��1�g��Y9{- %�?���|
�����g�xXN�\2/��f�8���Sb˜:х��1�J���o�~&��k(�/k����Ol��va8�Cu>��R��^V��~x� �7�x���5�/s���~�Z��p�{a��B���
-�ɺ������.VѬ�|p���~F�W�c���2H���V�)ń��j�_s���P~E�������|�0�A޺Ժ\70ś��u�����V��M�J���^wa��H"����&Y\7��M�/�	��mf˹��z1s��3G��ç���h��8_1}Tt+>��
Y���LGy`�
�_p<����W���*}ߺ^��%�AR��	����#�P���\���y뜄�v�;�X�E��>, ?���Vi�|D��M�7�kT@I6���|�Ըσe�oӁ���_�]$�oD�0�(e^����[�ዏ=��W�ɒ�)����H�h���hУ�ý�Ig�Hh�N��t�/3�)���� ;��uIG<ބ3��[Ha5Т!n�7��a��^����Y�G�7~�N	u�N���'�)��<%}i�0��D8m�l5���;:PϺ�^�v	����"̋t�ABe���L���B{Dv8�rk_J�4�#�0��&I����菋N�Ss���?#E�Ќ�	��N�q���s��z�v%[�;��bp�n>)�a��)�N��2�[8I�lL#9`%q�S.Ԗc�׷�Hb��e�(���#�+��?֢ȱ��x!�X�6*����t���5����v4���Kr4<�IlԄ Hʆ�!~�.��Ҋ6"�,P��	�����z�{×~$���@:,�Ӷ��t��=n��~7V/�7����������k!	���|e�s�?V}��x32�8��M6���9/���}-�/��Ca�����qY�����*�x#���h�FI�t�CԲF"���F��k�ԛ��j�ZL[�:�ڔ2�!v�1�QR/~��n��r�	��2��h�W��K�,k`H�@�&�	P�K$�W��4�I`���c��H���6?t�5+賥���9f'����w:����r�I[�H��M ��O����j��_dŐ���)�蟅��B*�xT�b�8:�+%RWj`I�I��Q��8+�{�V�Sp�Nt.��m�iq�������/�f<X����R?��0���mk��U��̂��ۛ��Nm������e�(�^ǨAR��9��Y.�B7m�����ˑ���n�G�a�u������M�R_P/�7���	�s?�~6�L�%!���G���� ��!��蕑�m�+�/���;,�\d'�vE���[\a+��� ����u�'x~R��I.�����&=�N��z�vmxtY�բT�rږ�CH��8ԖfQ\��n���; �D�Blݿ�Ȧh�������$J;5�`�PB�A=7��y��	ONp{5�ʢ��d<a���|86
4����Y����6q��5?K����Җ�f��eWƿտ��Л]�Ȩ��P�q��sl��o;zN�a�D��-ئ1^�(뿬v�eR�Kخ�;��a��K�*���L�����{�q��*�R��ݓ"�U�[u�U�,-�����,Tz��t�l|��t`����?n�N�wQ�|������q(��D�iU�h�p���.��B���KD�����(���Q���!�Q�kT�gTU�Ǚ����n�I�Ę�Rq>L�g���GF	�ss�!�ɷt��G5�ku���T+1�Y,
�GM���Ii˫�x����\�O%�t^5XSC��Ka7@�	��]w0��݅��9�N"ooB�v]S>���%ߧ|�,�����R���޻��*�ŢgZ(T5�O\ȼ�]p�J������	1�����0��\"�n�!�3��-�l0��R"��]�z���lKڟ��L6�9����QF��V�o����ܷ_5er uEs�������8mcxӆ&���#Q��+���B}^Ηtw߶��{��bO�0XS�^�OO���oH�$�6�\���v��W�!
�c��|ˮ'�����'5M
��&}H�2�-�043�ΨT�1--n��^��>l)lC��h�����X�&z����L�����d��+̤n�^b h�cډE�	|�
�F}f������SGW˹�<v��+��rԑ֖�ۘ�`{�t*p���~�Yɼ�-u���V�3F�{Fݾ�=�����ȡ�uM�O�,E��5Q�(�=����Yp��F@V.�3n�M/ �*C�$,s�ir2���r�c���H���,MK1%ݔ4֙����LkL�=��jm�[R�É��e��$��m_7�=��)f\`���������{{|kKn�R�6I%�L�8L)H� ��c�ц���*D5m}�HOV��jĔ��E�*�ݛ%K��rT�P����ꀫ�MZO�$�pJ�}~|vrC����깝��	���ۆ��M��u+�J��@
ֈ	�Ѱ��C����T�)�x)t��۝���p˞yx@
W"�ou�3o\/��Y�����T�6;W�#�Z�������91�(����2�*�c��c^LD��.y��+2�v�)�������	���u�&s(��O��e ���5��Y���=�Lo��{$o��O���OMW�\e���׸CGrF���(�DY�����ϻ��I7,�T~��6��o���PSu�����#6'������}2)ML\�O]��Hk����?d��u�!j��9wk���w�i�O/O�_���x@%0\rz�)��/�{�r�K��_9�M%���E8�w�r��Q�^K���u�JP�0�*����wWo����-]��G���TSaǧ��i�� @��Z��_��r��^N�w�b�>�d:�����OoC|�I��~��f���~$dQ��9׷�6��ve�!6��w�WyM�5��S�����I����W��[;Vt�q`a�4�ob����!4¤Qb?l�ʞ:Q�1��:k�g�E�:n��#C
�b�c�� ͐�g��@��#������7�+F����!�n�Z��.T�E�&̩
��9�������͆�r�b]�������$�@l�Ҿ���]F;���43%e A��Z�ߠ���Қ��r����Rݭ(�����.n�@��-�̕��`ˇ}���u\�ߧ&*Tk2��p�����Ɓ[j
F�u�9����0���^�^�y5�4=]�S\O��K�
�C`��S�g�:���J��>���3=��Jі���+gF��.�;VJ���Hl,�m8 |V��e:\Rw��6�ռ��x�X�_�"���@��S�t��XG_x��Zk�F��E��l%󶓌r@a�cË*����>R@����So$���<��i�����&�ML~�+�%%%�]�n� G�$�'	A�p[��c��%Z!�B.�Ȩq-���r!���m���ST��ׂ����v�	Ew�89TR���[��L����؝�Wq��P�B/䪁�+�"U�n�j�K�/�gM��͋��x�5}1�����l�G���nh�LTX��\fI���'9w|U�Ψ�~Y�'�;?s]��}O6�/=����Lj+�"8n���!v��`m<W%W��J�d�ذ�pA���9G�7`�=Oq��v�Vo#�y�\(]s��b�h͜B�c��iT��+⊁ 5Ʉ�l-�����������m����16�"q��cJ0��q��[��DnY�#$���T�g��SK�����xE���]���S+~4��;H��#���R�+.h�c\bz$��cc��8`����'�����[�B�R���$b�4��Ή��x��Bh�#5�	�e"� �k��Ґ+���P���>�~�>|��`��!]�I��Q��\��,��_^u����Vo�JM������� ޴�B1	�w@�"� ������m��T.�k���b�ԩ���؃�o�-���/�x��x@Q�%�6�����YrH�N�g$���?��Zk� ��l��N�|vTƢ>ߠՁ��N��y+甇[ ��-�+�ĶqS>&�h�ɾ���j]���mz|}0�n�
��*�_�S�!��K�&S��E�ZkK��E����	�Ϲ�E�)�;��퍸()���ǚ��N5~~ _��P��m��"�������kn�ʽ�j��2������0��Q�t���1=��%qNȂ��_�>���l?�8G4�=��]2����9���ǧ&�J�:�;�,,�s~���:�JX�x���H�ms>�j�3K+;+^��cs�T娶ވ��o(��р@��9T�T��^���Z,��\�_�W�I8�(�"~�?b0lu�<�bX�ء"�GV�8i"�2�VS҃�R�U�e�1��H��<�t���¬x� �MW��5>@�Y7{��g��J����ɂ݀����J��ślv��P��<	q�S�L9Neh�d]1�~h�Y@H�46L�0����`�|�n���=�uE:�D�W#
�*=���yD'����j"�����`>t�\��� d ʖ�˵z�b��%�=S�/(`�c�
i�Mo+Xl�I_��(���G���E�~�ӝ��G����hۅ���]��o��O7� _T������7X?d�},��ޔ+�k>D�B�L?j4��~�m7����F,.�1��(����[��������{�ZR<�W����`�ChÍd��IJ�d+{�>/��Y��f��^�$��j�n�/�Qȣ��I��x�fq�k�qC������)~�臯�q���q���!��ধdt,N2/(D#XDQ�0���,6�z��;uCg��s�����L�m{����c��jж��ӕTYLg�� 3�*@���k͑��E�������/���Sߵ)/����d�w�䢇U�N�Ec�YJ�h�X瓠��r��[[��F��{\C&(�`�S�#	�LS-����f��5���/��%G>h��z�\	H�f�5a
[��Q��N�ߎvT:/{��(3 ����� e��Yi[ ����8�}!��KT�L�i΃F��'��s����=u�����2��X �C`<�y����+˔E�
v��q�a����I	nG�dI,��G��Ę9-���<%I)��=���aOP���V6��j@���ND:i>��~7Q�����Fp;+gȊ�O#f�:O�j��ff��h����#P����[砞̥+񑡻�HC�9�S���r^+�]zE%\���3Z5��Y3��d�_�p�JQ3>$�`r N$�/m|ݢC-�����JU��}�<G,�����B��H�}�u���6]!�4�:+��h�(쑣(��[�:޾=k�����P+t\���5��_#���5�FN?e�u���Q�|���� ��JB��m`��8���=�����P#Z	JaU�I�qV8�l�8|�:��  U��sc�r�q���0Z֔*8d"*��ea�Et٢�e��<����ĬD׉�62�zm�_���a�w��>�6)����fj�k�#���e�/��>�EN�b-�~c���U�G�5�߭9PvDh+�E�!��~jcp��e�3�'gŸ�^#DF�BZ�M"�L��q�(%R>��+r�u�gJ�|}r�b8�#�ٷ� �\��`���^��.w����j�A�X0^T��_��3�Gt�����	��/��ۘ5_6ƅ�p��:�zk)���+�=�f�α�����o��&3��	�`ǋ$֣�}m���6 �.)�o�n"X�9��MY�D��9�C�b�;�DB��-���}`�N�6T�F��y�7O�_O�];8���9E��o��~q�R��PKİ*0;� ��N�Te]��?r�)��A.J�x�g�V� u�|��[�����wؙK��5O��MdT����+�.{E�Rb���Դ�L�e#��=�"��o�|���E�o��L��^׺���?I�s]#?�Zv6Bx<Ѐ���n�4�,�KH-Z�EJ�i2�V�E�=����13b��F�N��C�4x��ث��_��ٓG:7�<�x=�-� >!��<bS����|��'�&B
�: Q'�k<�K3�/���Y<�� ���"���8�pW��}�^F۾0b�h|~�ha�;.y�⣞�ڐWJS��U����Yu�)��{�Vr�����k�"�'����Rn/�C���^�8A��2��R���	���]��!
��}����̒iBd&��.}R��N
����]��w_0�g/�AgB08(�O�t����_F4�Wot���xp�&j4A"xp��k��b .�x4I(t:�#��am��~`c�3}b�Ĝ��8{��EHk�]��:���~b�@+C&�G����)���)�>Ot�'Eb��Ua��������.�y2�ˊ����O|�Kz������\�dy=;b����㇖��'&фȟ�gj#��R޶��z�t���N�Z�{��Q ����1^�{��p�g����ŉ��	�*U��`}��{�5�{ee��ʛ�D�(��Z;�W�>�!�o��)���!/��1�@R:4�����4)��T��EC��K����HU>z�k�a0��y`\G�_��7k\蠩�
�J8~�H���;#E�5ք��F{НWs�w�_���*�ޏ�< �Lq6���#�m>�xM�H�רۊ2;�"��X��$��;߶�`h^h�`��xk �ߩ:l�w��,�.{��_ó9<�;��{����z�c������n���xN��4���n��F����1C�ǻ���~(��T��`rc[<nU��#*f���a6���2S������p��X6�����g�X�+�8�2��C�X��v�%(?�L;�����	�-��~��dJ�*�O�L���z�5Mc�\�Qqb��WA�;����aZ�!���鏌���A	s�x�;�Al����ďYMGmh�G��� b�,cs�����6D�`Ċ�DL/��5��#,bˮ&R�Sp��NY"�'����S dɐWG�s謕�"�z �ˮ[��;���.��[@���D���!��=��C��#�KVCu����$��x8��u����<��8����LXt��n\��o��\�vS�y�ms,i k�~K��N\�ʫ�(��W~�S��?;�9[|��]�T��v"��~I%J� �u�������mՠ�,G���\,���PS���p����i�=�o���%�A +���H�OVa&@��82߀�>�����DU+s�]� \#��	<��Kܶk�����������ǋp\�X��a ҲPۭ ��w�l�pPɶ��ql�$v()5`B��P���p:�\�P58� {M@���gĠq���q��-D��j���Y��plP�������ٿf���`���v��2*�u�c���npl�~��r�h�?�k��W6�T�pi�y���Bl��l��U|����DI�i4N�z �E��c�p����"y*$�[J�	��Gkb�n�N ��{�j�hU�z�Ϥ����"9���}���<���s=���D�)�3�-���Ag� ڨ\���Yɫ}�:����S�}P�\���G�m�L��9cyu1ĉ��F4�k��`�,?�N��?ga��#W�'�H�0�F�.�Q�;zd4�k(M�d'�0_��Ԓ�CvP�iM�Q���k�9����'��Վ��j�="���t���YA�;Ȫ"��vU�ٯKp��(�LGi�{�3��U�ܙ�����Q[i�.�7.ߔ�#ٹ�)��FP���Av�����iL���&�wx��%S�R4�P���D��`hۯ�x����,'z@S�t�C��_�S�Н��&�PM̂TC�m�C	�-�8ɍkpS�c_����F�kɃ�?�~p�n�W�Q�	�&�J��O��$�H��I��6#	��^���NX�=ȕ�7+Y���?E���@MH��]S���ׅ@`H���F��'_�_@:�uL�M���}����<H8������z�mߟ��lo�s���jX�i�μ*<o� �Ta*|E��P�Q�?�c�6������r�l�������8҇-5_H�^�B��;�z�59�*���ZS=���"a^6V��$ n������m!�uEe�����A��S�*�-4��.���ҭb�ٗ/}�C�|�hc2�Y�&f	q٪W���I�r|%1�}��E%{�����S�[��[�8w�b�A'	(���H�Ң���S��C�A ���i.��.*��.d�zãQ�$���7�������Cz4Q��|y�:ϗ����լ1[���{�r�����a� A��I��N�I��"!([t�B�kg�$ ���"3&`;s�1�?�^�m��|����V�n?�#}����������r�>rH�- E&��71Ys����FG�8��";��ai�����
���y��r4MU�wHݬ�?B�� /~��}7J�BA@�y����0%	�k��eIp���ߩbs ƫ'1a�waKU-�m��&�Y���!@������Y(�'-^�5���`�H¼��2�߉���.���yܗ�R�e�?�MJ��밴|N��TDpr<����B��Bϒ�R8	ň)|K�/�����%wYX��|�pM�����)�F�-V3XЀ�`����'N���#� G-�i�D넕d�l�e�����)�奘{O��\nv��%RC�N�o7
#����< ��m�j_��/=WM* �W�A��}�,�j�V`����Ʊ�6b:9�n�q=^ǲIaI��j�jG�T���(��a����͡]�x�C��?��&-���=���m3�K `j�"T^b�	� ��gCI8V�+��Ɓ���^D1��ValOv��'�ߵ?61;�\������I\�"���&�^���H��r�����M8���郘�G�q]������'E��5�+2FK(���8I�Ձa��g�/;e$��#EiWl�r�Æ����px~��T�(6�*e����7�E�^`:O�k;���^2�w�NK%��Z�;�`/��i���1������ VT��\P��m?F�9�l�{40��P�����Ke�����K�����y÷��z)�%o�����+��x���=j�!7��p��ö��x��{����$�8n��86ĻS�R��fh����)��xKY���j�\���0����6hZQ��M�L���m70u��R-��6)���A�.�ҩj��^ -b��j�͡�������Y�m��ߨP���fB���bK��V7�b�+葇��O�J��U'����}�h�L��aF����+�nO]�{(/��	�k.�Ӯ#pҁ�U nъ�#��<E��\�ť���-��Jה^c)���EDx�!N�]#�b��C]fwL@JM�=��k9�(�%�o�>R��u|���F3]0��w�x|�z�w��..��cj#;W�ˢK���S��0y��T�zo������%��:RNyZ���m9	�]����uu��ּ�e�4��J+������4�h�EH�����B"1U���!t3dF-����^%?�RH~
�/�=x���l`�#�>r<����Kϗ�ѻ#_#���A�= ����G����I*._͡��\��K澌��k=o=Tv�e��=@F4g=EI���cjoE	�S�@�`)*�+A �Q�a	/Dwc��l(A̤2���e^����H	���ūm�Z���3�������2;H�u?��5�J�w���z�&�`�9���)&�3�'03�Y�ُ���˛n��<�%�bl�R`fid~�.ȅܞ�b���}�bl�:1�)p]�=+X����)�8�g��b �J��|}�\mS�#�J*=�G���-�M8`U���r��i�-!�]�	�4W�OEU��-L�}L�'�5���JO-�CW�=�慠"=)Do���{�-Z�O�9Ӯ&�J�kf}�̐���0y܌}��7@*�%���R�K��h;ךVV��＀�/��G�o�O��д���/���ܵ �Z����d0 �6l:���#3m�w-��o���+~� �VR0֓�F�oGV����VQ��F��Ǘ�;��߇��W��i	5����a��x��9������`E�u�§Uw�nԡ-3��sȉ�R���c��9�.�Da�p�E��+9xƐu��b��V� ���i�J�A�Wl��jE{�Ҟ�r,qD8cJ���F��t� �:�E�����|��ARU�)v�&���w���xY���A^��!گ2�/���	U���@z��(xmy��5�>�`�i����S7��k�5�Wx%z�>����?��sY���nKai�\󴈆��-}��'���R"�[ B=��%QY�_y� zԴk J����0m��4�ļPޠ<�XقmӮ�q3\᪺�C�|�rI�'mp0~�w�o©$����Aٰ�$U��2}�>aOG����׳_#�!�+�@�=
�� ,u(�^�c
�Bz��J��e.	ņ�+�x���t�g~�+�����n�]Qq%�CNZ�x��,�8ٛ���~���a�Z�����s�� l��:��V�4�BX[IJMph�MO�?���ɒMf 1X2&�S��?�5�p���% #b��9_[�
�01��	�:���������7�*�e�?�v��.F~��C�Ph描�2Bp\�h� U[�⣼��)E(��>L�2��t�g.)�t�泌݀�HM�W����s%
�(˫fQ��Ez�
^��&��v�����i>����C�k�5�%Z)f���>�&�n��H������3�'��VVJ)3%���R�̍/y.<$�����:�,������S��-��������W7 \�ܯ����.\�~���r,�9�̪�fw��n*�M�e��O\���uk��q�'oYqt_�F1��߱7�_���*U\���h�T^=.��N��;sY�T���B��j��TL,(�j��8��y޹��t!d����]PGUx� ;ǚ.:��K:)���D�}�r�8�$�,�B�u��
#p�
/�0ܯ^9wh%����Gx���)w9��<ag�/���2�3+�_���@�;'���\҃�т����-W�=�07�:~���o���"l����o�s���GF'�7U/��v�<.Ԃ1��@k��} Y��KE��ί[�Ҫd�ըkj��U�>�@�B�d���M���	�YCjNͪ�!Br��u�w�f[�7nŐ\䖞At�����"����Μ>a%�����;0����A��7��-|��D��tP�#�S}��u��T�2�R�{�s��H8_>�>�����Rz�Ȧ.O2�6 js:	�c�����e���l>�:�1���ŉ33�rz\�k���&H6�2���gH�L�vݦ�����!Cd,>A�A�����y�l�MK�0��İ!��E��q,��(�So�}���d�2�Pݥ��B-�ߐ���[�̫���Ӈ��%Jm���[�$�2F�w��ţ�_�k�1��UUe�I�>[�!M�H{5[3h���K�'�D m��:�m� �m��^�F��-����4��Nŏ�P6j���G�ܟ��q�՛l�N�^�Υ#�k˸f��l�Q�w�������R�˯��
��K�٫���@�����=w�	��1r޻�@����q(t��)�oC=i��&�Eτ�PAC����ހ+��"��}&\���[��nO�\=����ײ82E���y�k����7��B���Yt�scNO�O	�"������7�+"����ƃ����:{��w�����aoW
X��M�%C���W�xN�"p�cQ��^J�e2�-�p#<	�O��_Pܿ���3T̷m������[m�v����{<͗�����-��ENH��>�#N��Q(�!�� �#��x�S�*�H=��awW�����{n����=��T��W����JXX�܇���>~j��a���$�o����(��A�:�ݔ)�4�zC�cUȮC��]�����賂�K0�!wG9������aB�1�
P^3\Ti��$Qm��g�.��&3K���~�#�X�w���;��'~VC���)t�i�3�4��������t��������P�|p��_�ԩ!�D�2���s�d@��i[M',㮲�o���J�h�JUF
��3�US�@���Y�TK�p^��.�IMjx8� �A�P������t�YF/���7潄�g�vx��h�=A���E���ܷƷ�q��j��2dTC����
f��j	v7ݽ�9���񷽇y�S��m4�Qܦ�d�f�-<$��qso��H�E������m��\�L%�x�Sh��)�J�7m�9mH�� c2pY-7�ڥ3����{�L���|U��k��1����72��/Ȯ�r.�'�6��S�:c%��\o�=��ބ�Ŏq�C�U�y�?�2�F�y��3���HA�0o��b��9��9nC�����H:�А������li�cS.�SI>��ʃea��~����,�g���e�c��X�R�o����0A��S�~)b��==A�%+��D���B
��;�r܉�p����Ag���Bێ7܍�[�^Z_�B� ��˞��?g�: lo��+<>���`�\V{?5��ɇV��L�_��|g�˂�3aKS���fm�tv�p������uοA�!J�>:�������vj��qc�+�u��E���kCX�YP�j�`�
�7�tpyϚ���ǉw��O��k�_D�Q�m�O���7ڎ�����k�B�_�a7��e*���B§wm��},Α���Ԯa�G��63���ܺ��1A�S��^��*;���i�_�}�^���o��~�iA��Cn�f{t��
���^�rE{�<.�����ɋ�X�<�T�E=�"N�cJ��$�Z�i�[�G(6���R��t��r�w�n� Eo������f��;���V��p���f�\!m�A����ݽ�&.s�&Mgh���R����0��n��a��E;^�|"�p�5��F�7�nϧCj	�B�X�I�<F��ټ��M�д��2-A�r�����H���j���2�q�2E��8��1�K���}%W^��x��9Fu�\�,R�\o_���
�q%�ET��[ r<�`��0�
�vc�M�'��da��0�"���6Og��<F)�rV��Xa���a�z���p&J;��w�6�j�e��zO�h��l����w����%`_bߑ!�l��GN�k��p�U�r�e�؟���b�^0W�d��C�wU�:g�p�ǘP߭�"j_�J���ZE���M��GG�F��A�zga�S�A '�c��b>t�e� �m���t_�D��H����V����C�,��� �%���	�P�,�~�����)�E���oe�cTե�lGk�֨=�������*;�������D�\����ײ���i{8a��}Ę��2pad�{����2ƛ<����䕶�����;���6��|����5��c�2��PD:*��l�!��i_7Rq}u�׀�)P��>��\+��_|f`�a��9���c&��`]����|ݐ�~��-gG�:�?r�k�"��W�d���v�!|��Ds���}	��K�	�M��K֛�yNʧ�:L��^@N����*�26m�l��S�۶�B�W��@�8�Lu]3>̟�Z�-}p���I*�M�^����㵄6}tOd���/M�q�;i�6ά���b�a��%��0�"���˩�;���!&���+��MNb�Y�BJ`W��\��_��d`�08_�����8�[Ƌ�
r���J$�hވ�)��D���z�d��4L��c���m��mҲY� 6�a��>zU�TԚG|��<c��3_mZˎ�w [`68���~hƯL�^Tׁ��c"%�>����<g6 ����G&����}V�rTw;�ɎW*���2�H����%��7�?ϗ�B:��}":�:�/45�HA�\d]W[jzQ����>c"��d������x�����ue��OY5�BP�_�&�j���H`�r��o�ۛ�0��6�5�x�w�GvQ�h��0��չ��d�Պ�0��^`�	8��:m	,�ע�z01��r��q%7!n,"���m��2���?j��.���n;�r���P*锛���Mt�GP�[����9���$�ҡ�܋-!,�,2o���_W�����nDF����;H{��{�׈3M�-q����boJ��Ԅ���T���Z>�gر��{V�J�i��9.���:�# $= R]W�\;̗{T�9f��
����oM����9S��������Ʈ`���)����M�Ѫ��z���5�uL������;�O><N��1��$���{�6p��O�RN�G?o[�����A1�3I�N����PGb������^OV��mx�)��/���D�z?����mdn"P`F��*�0�D!�]��-�WfQ�s�5۾T�G���:88,�G�(����v��WL�+���'���=���?�<�3$ޠ
�SO�\LxG�[�'
�����|�s��T��x_�0���<I#��s͛��p	���y�y
�s
@�4��8���W��>��of���ǝ
�uK&3'��>Ot�"��%c�׊���m��L-�2��b��)MJ�F!v��FA����_Y���Ү�h��7I�d-�*5�ѬK�?��:�{#d�Q㉼�`y|c%R�v��q��%��,@��5x��e���؆b�'yü�������I~�C7◿� �L4�U�4��z�PF:"E�� [���ꢃv�����4��˙|8�!"s#����2$$mE���Ժ�VRW�p�{��d�K�ǇP�j^���oc�������e��,4�.�&�dX����(�D/Em�z�P���ґw��b�4�(�d�����8�y�����;�Il��ۣ;��~�8�z�tq0I8R����EAG��\@�Yd&W��OܩU� F>S����.inF-ǘ�0<ϴ��8��zX0
O��E>ډ#_�E2��0%=�My��f����u�TM䛛���