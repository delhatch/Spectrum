��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J>E��
�L\�īi�p�H7ȥ�g��D��W��(����'�yh������a7���	�'U�b� zv��_�i���y�ǅ7����e�4���%GJ�1q�>�����7��-�7ig4n�^pQ*,n�	��q�K���w/(ʞ"r�����F��g��&sµc,�Eއ߼�R�ߖ?��첎���~+������߾� �\�3DC��g2�6�J�ڍ6Tج&����6��s�v:
k��-���]����g>r�Q̾"�����ǫ����>Oxv�ƫ����ʄ���o=pI��u���XZ~�\H�p"�ɱ��a=�2��-}	4�����j������r�j����31��i��폡������dJ���-m]���Lo03�KX�O�B�Ǒ%ӥ.	룥��6�Dl9�/��t#:C���&X��w�_�pLS:�9�������7�1��q�NZsp<�������M���ޖ(��>�	C?�_M��u���x)�Y��2Z)�����Uݫ_ݸ�JA�!��.��ZR��ږ�fգ�;�82�T����90�^o_(R�j��HOj��E`�8�'�ϥ)e���T��!��R���uE���M�N�/�|ۄ��F~�(FV�	3\P�b�K	���0S�I��vi.<��4e�P@�/�g�Q�m�����rTS~��B5��B�O�)W"({�p
#�/�M~I��IY�XS�����W(��U�A��J�W�r�A��i��q��z���� �'�3��7S�vp �\!��k#�+�#�uZ<U���a*Ǔ����R�� Mփ�y�I��p�C�>�_��z}	W�,86VB�1Q?P�d�?�OT�7��������if~�M��2 vo����Q���|p��	�v����}�E��a���=n���RBT�]ִ�����dk��ڲs�Dl�R�h�^�<*��ţ��i��rTF3�#�"3�C�ԂX�r	l�]m�=	���&l���s�+�$zN�L�f#�~��+È>-YfB1V�a�{rJdC�ŀb�:|u%�dBvB���mIN�w̯y�����q�16d*���E���zE������$����I�IW�W]�)˻���\��a�L����QP���Rf�[D�t;c55H%;DD?�������O�A���$a�e���耪��Q��SG)C���X�y'��$YGL����ڞ��XS�V��h�����X�j� O�7��77U�:F���q:��l�=U�g����^���7�<�CV�ì�o/f������˧[�����Ml�������'p���7$Y�5�]�����q�^��3���_9!��GhXlb�p�lEg�Z	��
jǢ�$��K�Q��J#��{�Gb�ݞ�{�z�B� �b��/{���p�О#Y��_2Q\K�s��<)m��r���yU'�O򘅵� ����7�b|����~�H�� $����+�f����OphV�iO'�1���!���Ȣ�FK�к���.�0o�RF�����Zbs���e�|�B^8D7��������&�K.�5*WdU�X��c��&����]x�!k�^lD�k�QD	3}�.k�������D�	�A���D	@�p�jA�F�}.`�����
���X;��ˇ�(��n�[�(6�D�P��W�},�F<7�_�3O�<Nd�z�����<RX�0WI���M��J;���8�Έ�67��ؼ��J��7�Sp�����n��B��g
K����-�rM�;�?�_{�8$����zu=6іq|L��ŉ�j�_B5��M���ni�'%Z��9�m�{T�84H�Be��E}��\�#"���q�Rz���l>U��>��?���}I7�B��Hl����Y�!�*l6�|R+�����$ѷ�\;E9�j���om(�����QQI���8�=�jf�]g��ApB)���뾓[AO0�o���.{��~H����d'D��-~�H�4��G�l�EE���{��<P�oi䭙�^� !���&���9�K	��"F>~���=Y�m	w�(q��@��w�����8oz�����-Y��T���خ�E(w��̬������%x���Y���'���S2p+�7Xi�Z���������R�n�? ��*5aDGH��0�:<�V�C9�?
�������$=�LV�?t4�( ���r�p!J��$Z=M1��T�e)��h3�X,- A�y?���lOtnN�lW̉OJ`\W'�6U9ahk;�:��`x���N������G�މ4��L�}*3�)Ӭ�����Y�>ot�u��9b��M/?I`��=֪��'��=�$J,����v��]��`m7EF���ؠ��K��5#�T�[�w.h\[c|ņ�r��lu=��!��0�"R��o~���b� ���.�����d���ʨJ��h2�A�4��i ��1��*_pL�OR�[1>'rt���6�i�X���w0{�0�v�^����G��.���^so���D�h���k0H�bղ'����5h�ɳ"��;�p:�\���7m�6j>��M��G��� `% �	N>���z�@��J2��dYF]��g��ݣ�{u��7E�k��Rn��X;u�<���