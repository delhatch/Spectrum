��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z����#M��Ӄ0���MD*F�L�>�t?<$��"��@�V�"q}�s��d��zD B�i�`��e��bƄ42f`9c��TTV{��d�!c��>�m>���b��z�#x�ĺ�B
���/���u��!���~�_�cti�n9Wwu~6g�Oɍ=��m����,9��(��H������zM���$_�?a��)d�%	��s�*Y��!u͔y(��dD�?�2�| _y??�L�/��Y�3�\Yg�Q$�닭i>5� �K4�E�=�a�λ��5�}��.Ꜻ���<�f\^%�ݫ�-�:dq�/���[?�!���.�	3���Eb3��	PamV��|(c�*Th��u4��]�2~��]�K�Z�E��_�L_��8�ϲ,8�b7Ѱ����r�)#,_���s��/�Y�N׳%��Q�!���`�<�C}������ċ�5$��8Y( 
���Z|2/��&�ȷ���sQ����q0Z��+����c�q���[�5l[*����v?7�=lMZ�eרX�oaL��S��N�P�\VJ��1!�]����������k�i��v��wڥby��Q���Ɋ�A0�x�����K��C�w�\�M�H�FRt�������`��ŝ- '(Ň�y}�v��z�0���
+�Si��B���3���R%�,��dfOE�GMœ��a�XV����%��#��݅�WN��̴˥[�Q��&�`&Ӿ�;t��R?b��YY����[	�pK�rzK�"��[H��%pZ*b�ƹ˽��b���ڟ��H�݅�jz5"�����l{��B�G�O|�F�2N~c�Dy�9�����n�Nj�Z��M<��,����[�+��M�9�ܑ�e�z�>��`��w���D���5�=^�����ǲ�k�p��Wk%�����3�{�Kvܰɛ�����0[P�OUQ	S�48ٹvRj�����Lo��Gf�#\�/��ϣX&�ª
�yJk�����5���L�]=_+�����a�^�}^w���3�*���E��Ҽ���?�e��&U��N#��;�J��-���b�m����GT�WE"@x��ޑ�E��Z�֮��r�/����W�Ԑ)#k9�q�R�F�u���F~J�~�'�u�AR؀��BIIF�����W�.6�h�����t�DVF�R{��%<�rnN�'�I�7�R�"��o����s����i��9��I[�/��m��F1���Y��3dB!^Awn8�I�����? ���C����!ڵb���z����2��?`��_��Uӟ�;x"<m(y�x]�0Vk�A7Eq���x6��z��o*A;��j?�/�	�9 ��U��
=,�X+��~���w�'�7�֋�����:�]�Ս�D�C�A���<�gT�}�@|@j����P�z0̃����D�
�kjB�{P��5Kxm���J�����.�3��_�^A�F�P��������c�� �jY��;�'�����0�\|q&R4�	,�ٞ7���fW	���J�K-ܐ����-��:ፓ��ؾ/�>�j��X�����۽�S�B�_pl��Q�7f$d,��D��2����+��u ���>�f!T3R�"wv,�aA�E���^=�%����ZV?yQ�	߬݀B���m��̃s����J��5B1*���\֭�8!�h�J:%��j�P�`*_{
L��C�t�rS����s���n�[��?LA�*;�;1���V.���;�+F����+�K�q#z.�����?���^���1h���ž��?�Ӡ9I��P�@	�J�J�7��5��:#����~d5�����G�TDs���ާ�$�6���'�CY�H�A�K�N ���Sؓ�M.�p�:�đ{��#�� ݔ�q��4)+;�O"�~1K>�,xϾP�����/J��/�8�#��N��^�6��V��g��F���<k��d���B�����}�|Ϩ��J��[Fs��hz	��Q���v�fa|1
�h��wNL��N�j��yׇ�!>7��gLv3�I�xp�����6d06��c�Sa)W-г��og�f���%%ݙ3����kl����m�;8�ޚ�X.�����-ؓO��>鼆V����kc$�JO���.o���$O4GF��'v!���f9�b�Vu�8B���S^�8������Y�� �tf����R܁�!�>�o�z��r&tȳ7(���U�A���7��Z��R�BX��z%���Y��%_4�=&Kc�}�G��&��_}w��E���mn�nZ�=t �}h:�V�<"R�9����1�P1ۈ�3��H��/���6kq���d� ��Qǰ5o��P��Xp�ߏ n���vWm�+�=�C�5�%T�N�m�'bz�:Ȼq
W©+[V&69����i}������~��i�h ]1m�c�Q�V��i���7�f\[��3�+m�b�
�r�CHF3V���<,Ђg�E��/��Gca�E�U4>C�1ރ�a��G����J��*��"vMt��77�.L�k3�#�_lI��G�Y�x��"�|�$]�*\�t`�M��T���:c@D�k���F�J9d�P$���"=���6KRV́�TV��ex�o�k̰�G�+q����p66߲�rL�j�$�аoH�S��� T&��I_F��L���㞮��1�g�·��Vy8�S~�(�k�%Y���I?��qgG$p�d(��_J^Z\���|H%�}ܗ>we0��@���w>���=׀(78��T�T���'� ��ͩ�Y�%��O#���&"7�#��s�� 5^iZN�9��9w!h�0�;.ԧ���[���܉z���X@Ɋ���L5'y��M�� �q��J\Nf�~��1����|]rNx�ü0�ų.��^EB��E�����Ċ��	��k�(@�/�ݓ�G���V�mg���1�]�k�Qk�+�*b*�A⎴ >bR�h�x7�1i�.co�)?k.PAp�t��o�g�d��0�^Pc|iVb㢠�+�m�u6��<V��L��P1�e#���4��0�s걑��c�aV>����?�Ӕ���D��'�y`IG�ε�4��� �a��n��X8�R��dO�yW��+%\��~d�*�dҒ���~&pvMsI�k�>�C���׃7�Oc�nX� ��J�%N��C��d��(�,���W�>߸�t��D%���Ɇ�Q/<�RfH%�pE���p��8�<E���M�w��p�-�f��xJ�^���#�|Poe�,�n*}�ǚ���wC��wSk�(�U�ϯ���O�) scTX����Rv�m���ϧohLBJ�g��Jϙ��،�4 �(F�Jq��.��*��%��Di�S�����;�F�3]�Zs����̳����s��j V��"��hR��Ҿp
�Q}���\��x�>�<W�N?�Ƿ������=JjU��T-/m�5���F<ǝB���N�p�wB�JQIp)�;��m;�Q�x��F������!�g�ѕ�{g=OhXXִ�ⅇ�S16��������Z�iN!����.jI.���E����:��G���tj�!.3NF��W�e��/��Z��+�w��0��L��!��qK���ǜ��v���)aMn_#���ƁO� {b�rkƆ|�h>�M�h(��L@M���7!1����8	؊jHS������0���EM+ˇ@��r���h[La�<���60���gN欲��b��E�_��^C��ĴY��C�@Π@�k�;��h,M��G��U3� B���S�6?ݦd���xa����qڰ��dĘ�dO��f�]�{����X|&���$��/��f����1������rKŸK�&��Vww���������ɒ��s8��L��K�e�3����K�ܗ/� ���+����z�-����9��7����)�ԟ&����ܦ'[�:���)l!��e�	�.
I�H�^��-���+��W��?A�^#S<>.�6��lfwo���O|'@H��R_� �y��@s+BzG]�e���l����C�jT~ܡ���83�s}��6�~/F� �2�/�}��]qg�}$a:�����ؑg�&��&�����[�do�ڋP��M��E#��%>w����̰ϡ�&a���Ⴣ]�P$I{t�\Z�@��l*ݻ��(��0����� weg�SF�q�'�*�o����r�a2L�]Z�ڎb���q�Y�f�+������}������J30�{<N_�*rvPQ�`�Ν`�h�{��+e��nC��Hm�?�u	���F~-��;�����c�P�݀��,��+�F�RW�=����%��HGEN
yt�����l��ֱ�b��.�A�,Z"�<�"�:5��H'���VE���MYĥ���W������h�U�Č�����\ͨO'�b�����w1�X�:/�!sNn��Z�_TԖJ��h��4�Jj%�n@\��� UL/��-��}N(����X=��2rq�ʬ`L��3��I�{ %F&��H%4:���PS9�ߡ���l%�Y��vK�%ѕ\"��撴|�߉1x�	B��>W�����s��h�9׌1)�pR�Q���+�#��#�'�Ҙ,�2�Gٞ�d�/�e6.���u�/6UjqUa��4l�	�v�\����T�tQ�����3���ޤƠ���s�8�L���5���m�])G��ِ�3ϋJ��W�L��� Md��#Ay�}Uȇ�u�������gNj�F�rJcH��<d��y�"�zWcd�$�k/Me[fp�K�\nm�G��|�Z��LE\�6i�/�q5���0�rP���a�i�=��ꅜ\[9ڕ�k��.�n�tQ���7'iph��/�kJe��<?��l���z^.ѽ"⢜���	�/�_�9�!�����ft����*vu�(�;PyA�hB�]��uMO��:�m�U�.�F>N�ܞ�<�L�3I��l~
�=
�h���;�~{G�(��#�ƿK*�A5�:��z��ʭ�	����<��(�BC&�L�IxP�7��7~눘m6�]D^?���\�;�DI��������M����K�ɍ&���j�;x\>Mk-"K�2�i���*'96{]di�I�7���B6m�5.�6�|^���L����`5 �g�u<�ݸ3�m���?j6�(�y���=E�V|Ҡ��5��AG#�+/���6m�W�}���]���B~Y��Z��1㠴7ÿ�'>r��3���́�����	=��-�i�����hyCF�b�$kz��%�4`��|�IH�y�?~��=��2q�` �������Ǽo��8�3%�j{��/��R:��
)���cM.��Z뵮(�g�����'�QY�����S�-+�0ۙrh���.:��/h_�!��6�͉Y�D1�O���G^�4�?P7���Е#���}���&�qMH���^�Г��:��*&������P7���2�3����Olcᝎ��*�3O
q�|���m�0��2��k�v�R�o���5�QUf��2����8x�2u��CyG�������]}L���4�n��Vf���MXW3Gx��xY银��`F�S'���x�ք���]Ө$���Ԭ30���M�zp��8��A�f<x,��3��y��%��/��;�
3���<�[�q�M|�7�����aw΋�f�
�\iΙczo P�ۢ�Q��D6��"q���1_24�����K�֐O���SE�?a��al�E|���>K� ��0΢y%�w񊥥�>��M���l[��§�~�'.B�1�TU�*��b9"��Q�F&��(>k�GVpό1w�Im�����5ILB��U �%e��VO�����1M��[�]CK�K#�qmX9�+:�W�g'��w��T��7c��Jj����O7�5�{:0�Sy!�@V�mbGGYq����2�S<}���t���'���a��#3R�v�!���<�vo2��q�ӱn�����c�{g�q@��J��B2��JЕ�]�ɓ���ނ�"ԡ�jŃ]NѲD��X ��S͍�RjIǑ���+Bz���pq�o�D����ǵXH�vr��Ϝq��å��E4��R&t/O�aa�/���ųvY�R���w�<n��R�GoPt?@[���{6�-��Bm��k������C�{�h��r��ڃ���X�Ff��/2��֖�-�z܈���dj&Kap���B�[;���h�1/ݓBu���0W��M��_B�����p��I$���������Z��m���hE@Ux!o.�̈́����RZ29������,R,�%]�	�	��%�[͔�G��Ӽ����xkq�uP�J�,)���4�eȌ��|	h��<����N�0�IC��M��£�ȝ:������>p�Qź9�j��2���F��v�)�m��RKt��A��J�'z<P�8G��0*A��^�o*�%�#Bd�=~�̽��$S�R�)�wJ���h�ֈ �P<�ǜ�]8���������l[����WP�k��Eg)nF�B��7�w��5Z_�Ɏ�M���%u�$&��S����S_ޒafy���u�K��bX  ��t/߫?�7� ���]opg�m�������♭�Ah�&�H��l��xjj�S� ��} ^$��3��;��IXf�!w����y�?@X���i�HƝy����$:����=�)Eԃ)��,��~-�DV1��bă��X�-ѐ�A1�zJ��3��1��S����dg�����p|s<�9T�!{�ٖZ�n$�NPF}t�r� 1�yŰ��F�BN���.�7+�y1���t7j�byB��f��I/���B���O�s�����q�7�c+=�~H8��H�|zm��Ǆ�9����G�a�Ɏm<�CZh�##��(-�Y�pAٗŧ�S�߷0���jKe������"�}Rl�RFV��w�z��ui��mT��&H�� {^Ns��p��F�rFQD6NqTY��ǆ�V�%�j!�G"�گ���t�]�xP�!ڽ6\��e�v&�9��W�'G�
F��O�X��U�W�`��A���~t�Ҝ�w,�T*��a�l���0DC��P���*Ԛ�M���о ��cW͎���0Y��h��v#���.�\OD�F���#�yǝHwV��{��/o~����sk��)���ݟ�CA*QP��~;���"7��u��X2[�I7����I�m�\�F�[@��>++ϡ��W%�����ц��^�V��\��q'��{�q��Rۇ_��%���s��j�'(�j���FD*Yy�J/i)��(,��$�P^Z�w�i(zS���GZ/��ɳ���l9^C�鐃��E�P��v��F3�)
��rs/;s��u��H��B�U��`���)�����:ѰvƗ�{��MP�S,�NN)}����E�'�7���H���Wx�ʿ=H���4��(���9U�%�n����_�%��Q����p4 J��:���T�& ���x.s�����n�����h.p@0�>z$��L�� �S�Fcz{��U��3�mvT��z��Le���X�u���o爜�s����~��xb�z�m����&z1=3F�F`y����!H���é�1��=�w���*�-8�+}�j�����-1�P��f�r��\;��}��Mۅ.@|Nn*�y�EE9�'��rσ\�ȝ�n�V���,m���Gj���@��tt��v��ç�㻀u��W	����"-�t�/�46q����#��=&�Z�\*8i��⩈/�p�;@��h)�LWě���A�ͅ�i�ڻ����-��*�k�Y�l'�L��カ��,&s��n�g�Tx۹(>o�chk��@�.o;�M�` �a�uWDi���V��Y�&�􌔩�`�$T��Ƞ㼌!J�$�L��m7�`Zi�֑��cŽi��7P3n��k_��.,���O��b�)r��@�[�� �b�Co�n���Љ�+�$�BX
�%N-4��S�\��� �^]���~��IV����X��Ɠu��G@������q�}�4���zm�f� W���ԯ���ڇ��2��y��k�g<V��u����`���h � �7�hp������+�	���4�~/��Ĥ�rw\v�u�_KBk� H֓�_M���8��ٹ��4�j�^4���T⺳��>��B�6���h�n��6�2��
�U���u�mQظ��|��9F�n��>`�-���%�$�oy �lܔT��.�}Sg�u9��\���)� |.o�i�	t�7��y�T���k*�rjv(��`DK!��d7���'�������O�q�� �p2�-O|�au˨3��QiV��#L�Gh$j6��\Bͳ��S�!�Մ3���4�bB�����Yy�3�y�tE>Lnl��	���y�,7z}|�ى �'��T���Ȣ+^�r�[��SX���N�2�_�o]��i��j�s}����y�>�1%Q���F���2���wWJ^�S&tt����? ��8���t)D]'m���i�7kP��*p0)g��qC�1MJ�!([�Y�&0�
��AQ��6|����Q�WܨИ=v��9��Dܖ��+��5]5��Tp���]nl\���"���5c�k|�S2��A�+e��l�)��ٓAk1�.rX�1��>{����8��:0ۑm>��� +7�4c��̢�#d��x-)nӎA­��¤N����A�%���`�*i���Ed4�Lx�;�ʡ�+�Q3���~"l?j��c_���ʓ4�<���fp�f��S�Tt�d�7�ו�#���A ��ľ"-^Y��]���x�!u ���l�5UṶSw4o�3�a��H��\����n�uہ��pn�A��C&
�V��J�������\q����bS�$YJ��y���3�h@���o�9���M��ǹa�&Y���q]�����l�O�|j�WK�`����ǌEgO���� �3���P=�-���B*Y���WP"f`�wv�dNFa��j)�TO2z�������_�" e`ʐ��	5��x��ߺ7��$9��ϯ���8^pS�V���H���*l�8����?�8�S�. =�٠��#��h���3cGN�?,"G0i'���7LhJX[���Ǝ���E^ _�v������l����3W��vzj�Ʋ������ӈ�D�_e�o�*�U���(pz¡�rZ-g��r�6P&���&f��x�s6
[H1J��O�)U&頞�g72i,`Q��Z�%�0��vn�ƍR��+�䳆���mD
~� ?��L�Vv����H2|�,8��{��4`[F�e�P��H��,�ȏ��:5.jalGg%�@9)���/d��UH�����ImsҊ��<x{�(��1�v@��]��P1-�=��Z�JߕVFhrb�S���$"�d��B������D�����L����m�(�DU,����R/��h;�N�0
��tו� �sUB��/�\,n������U����@��h��.>����{/���7�����M{�%��184D�f��F���ɶ(?u���F8���AY���>�[W#"��b���J:o���B]������T��F�Q(�QC}ʥQ�`�Fy��-�1�G�8���HR��tf~���R=f�#���?��y �<�0���ݼ�.�I�TgK��ޡ�xa�})���e�k)?�{m������H�h�vV�q{$�GBO�o��ұa>���@�VU֔��[�8�5����\"r7�o�����ۼN:�t�b44�,Ǒ��
p��w�F�^[qO�A٨�0�o+cKTa����'d��h QV0�f/��xp�}ٙpB�/gT��/O��ѮΕ;HxK�l\ ox�7z3q	@��¼}��;��4�)Cp�	^aR��V�^��������wo��JPS�fŬ�)	����f��K��ڻ�{�>y�<�Ә\Ѽ� =.3��/(׀���?o��`����r��q��r2$2ً���P��%p
��5lL�<����#\!z��+^XݍD_�� �EА!L��#H3��O�ۿ�+o}
�6w�ܕ5[`/���m��ENtT��R*Vg��!�Fc�~8(��e��w8��U^)X�����K��N�%ܲ�~�Y�"�hI�9�U}{7��t�6U�̳�K?�.]������?gHι,"٢Ȟ�+������x.W�6\����+��̪�'i���B�ˢ��*��<�� �D���ފ^4G�ƾ��;<Lg��F �t9�I/  ��{���P�XR���ǭ,τ�ATRO�/m����{���í?p�+��q�73����J�c�K�#�䠞�����ƍ��l��5��2Wif����Xm�`FR5�K�����Ɏ�`N�JO1�Y!3CF�\��ǜ䏉��z./�hwם+4 %MP�޴�ot�_;��[��;���j�a뜆8�0�0G���O���� 0�j����<TrՁu o|��2����l��w`Uxzg�S��RNi��U��.�ӗY��Q_]߂���'���bL��Y�]�wsъ9bkct7����q�~5�N}�N��fm	� f���;��Z"��īw�T���9�!v����ɦ�DJ�p��h旺�wa�L�u&'53�S��5�i���<6�9�j٤BǆW���u����6�0�YEbz�l��������T�@����x��s����Z~�|쵭x��"�����{�8 .V�{4���	�w#�_~� ��'�t=ۙh�J]:�/�Y!2X�-[�$�'̄E����U��|B�S-e�b�5�,��I(���!�&��Y&#�B�5m���6|M�rKmLw���U��&�@k��}�f}��)�ۥ^։{/j���WQTfz����{�`着�M{R��C4߅&|�n�Sf��(ld���)p��q.D��*	<�O��.����N[nf�HS:	��&�CT@���tO@�G�¬6��Ji�(���9��C�Q�#�Y���!�sfW=Pq�Jg�X�7��f�o�ÊT#�}W�X�kF�A��4Ľo�4��m*J
�E��.�ĳ
�qZ�\�9�'�:��/�A��$���l�9�����O˦R�|����Q����/��%�y�����g�?&���ԥ�2�w`+�/�؈<L�˂�� ��z_�k�����j+�F���,��F�vJI�)Fx��D�;��9z�G�����Lox
�xؖ,�5��'�L��J_��_|-C�	Y!��	e��ƫ�YR���tku�x���TCL;6^���!��oF~ňj:ę������q���9��yZN��\xF2@��2��D���Z��f���K��%�}�V��)�_���!eY*H��,�l�c��wy)�K3����Cۥ��2B&D/fnQ����TQE���u���68��O�%��sL�]}v�_�{�A�}�15bX��ⰱ��Q1
�H3��K�F�3H���-�*�j��γ%�/��~��8և&#d}4Ѣg�c�M<�g�0Ksg%?8����L��\��ȲT�7Y'�K5�Kq���W�I0i���.ֈ]7�H���	����D�X�H%u����Rȑo��z޺��底0�%�k�o����	'�br��/�]�j~SAo��g�3G�S�Pqz�$�d!�������FF&�s��(��0z/��~]3��㪃��e���E{�B��V���+�܇�ɬ��S��|S/wӉ	�'��7#�t˨�d)�O*9�
^����G�&5�bh��U��l̝�
��]��?4���f��:mE�y��m�x/Կ,�?�}�ɑ>*� > �A�A��h��m��d:>\J�f�yr�O��So�n�Fƭ#ή�b53��-�#)��#���U�R.6��[�n�^hs��&�c�=��C`J��Pg�������0�� � ��-)C�6�%�G>䰄��S&��ڱ/���?���3t�=2x���o��N9�s�g�
@�Ն�ƤKK��k���.O�,�1͂�����]�(����u����x�!�b����~����r`�[td^C8�ќA)7��%~��J�~Q����_Z�;�W̴�a']ػID	�D��� q����������^ K��@V��u���R�))���<͌��N��1YC2�A���n���j�����Oc�OF��Z_�{�K#=�濻�������a�F��tä���$O�;�����wO��4��ow��\�p���l�����/�p>����Hs�s�XN��{E�5=ɂ�I�d����Æ�x����J���V3V	N�H�E�2I�冨�a�?�g����>�J���Vf)M����������3�L���e��82��]{���"�ǔ9�����I�����]�S��p�ˌ��x�g�>��A�T�5��$�'k=I�LY��iW<�����I~c�,B_th9�n��0	�;<̣�;ěD>Ϭ�>��È�5p��`) �Β{�jnh��M���@����Mo�ɏb3
�9�>Id_Ը��%��"�}"����f|�N*A!��?eՒ��ꃉ�(Wڜ��T��+Xq"��3l: !��M��S$>iC*��#{<̗��f�z�XS#�*[�jKa���e�2ܠM�_	n��E�/�	MJs��w���X��旮��x���F�]#�8YN����}���۫����sR�I�x�ж_�H��J.w�5��y�^�2��� �"�|qX�3��R6.��9q�t�ۼV\�g���6*Ls�kV�Hd�~ǃ��<Lt�_����#�|����m�\8Ev�m=�G�W�sG�39If���l�~�t�eH�hZ���q�?~���ZS�}�2�8���'���i�:Jh�������=����>��+'�\��v�d�S��$����Iwp��ƒ�.�ˬ���/�f�y����j�#G��	D������t ����l�MW�u3�u�{9��閍8$;аL��u��׼��� oyN���3#7Ѣ)Z��__ઇ�e�]Ә T��>�(�&ʁm=i��x��f^*�%���v�� o�K��&\�Spn� �;��o������t�j����9�C�y@�L�;����ަ:[��+a[�=�-;�O�2��$�QW�w�w�8�Z���;8M,Fbע��!A�ƅ����'ͤ?8Me�\+H�/��p��U�M�`L�'������z�;2"K��`�=D@~������$���#s�DM���zW�ٻ(��J$Q'�pj"��t8h�����T	�,�aDO���F༇e���a$��GtqEG����w�N���x�W}S�J�����͡�������҂E�c���J Kn����3�{��C�(Λ`�ŧN���n	p(aU����-�v������ە��p� �Xm���c�u&����m������b)��N׼�&H�ZwAs���)S�33P�̆,�ȡϙ�k�S㦸��}%�(����Y�,ճ��}梿E���V��犔*,�.s��
]���1����T}z.�1^�R^C��۹�pw*�#�	�n3a���`hx���xƳ�� ��و±n��P�|�١�y�W`��Vޛ)~K�i��U�{��d��=[?6�{� �0$���:J@�!t­@�dWV@es<%J�t�f����8c����^Wz�&#'Dj	b�����t�>i���=Dq�������KZ~\�:@P6<F��u�v~�#���;�ǭ���+F�p9�/�B�7L���\�%���!��n����Ju+~^�9S�\��\�9D��&�?�&#č��9k
3��"e�I�o�>�+:�+1ǒ?l��k���Y[w�x0xa%� �3�Hs���y��J$abR�5a��M8�Z��?_�K�A�y=�������իcǑ@�
�ě������DTb��y�"��^��FuN]O���ɘ�iN5s�����\��"U��3�{�T��*�¯<K�3/��~�{_{"ayS�����Nx�Ԥ�۹ɟ
�(B�ᎎ�@�q��%��$G�ܲ���-2l|�\�����9�5F��	.�)4�J,erJ�+�#Nؐ}J�����=�]�_KW���E~���rh�ښ�#�`��
a_҅EQ�'1׉�#�P]dT�Ioe��1�͝H�������'��V�T�m�̼�G[�)�L����}�)m�']�S4ƻ�;�+��Z�3Z(�³E�0[ju�A�������6w��	���*}�{����Y:-N�1r�z�Tҕb�
Tq-r��9t�Ť����R�a��[������/�Q��<k�]w`)!�2�$��w�UZ��g4��"t9�6! :�ә�p�����D��+���\�n��\w)�F�Z�p�7�"�+�)qg������̊�fh7L.-û�aSfg7)�z�g�e1DI����*�Ρ��^7X���R^�DY�Ó�IzI!���%9ᐅTW��3�	���Q��J�(����_�ı�/�|�FD��}��9 ;>��\�DA �':rAE�C8�ȣ�@H��o��z��;��}��	���!.��[�9l{�#�SݚV�����'��>��u�b��#���Њ�k��>]��]6�f@���߮������x\<9q������t����[�oE|R޹��y!VwY�C���t��,{���Z���w�����'���Gj�B�"y<���S��˲��h/^6�D��}5��J���*�f$��?NWO��~Nn����N9Dsi� }���j���iܡO���,ʚ�\���,���S��֤51��`��BMlB���Z5=�QO�iG2����Gk�TO�V�N�����w�LTT��c�rR繁�J���<�)1H���B�w¹�f��)h>x��,r�X;Y��:{�R��10�_���	6�H+�)�Z�\b�4�Ad*)g�s�%A܇˾8<_v�î�������?@>�W�N��i+Ns�b�BG����ۂ�j ����;(Ƿ�c,�(tZ��P꧌%�?v���A�˯f����&r��
�eU��H�Ǯ��w�I��s�r����������ʳ��-, F�=�S�3�=F^b��M@�3؟��h�M���%W�,��axI�ɘ��}��W�
�[.Y��o�eO�k6C�"%@9$��iݭ������%c���C��d�9t*��[�'�`��-��suj~0�\W�b�-�z���z��ױ5�Q�K]��g�zkDኟ�j �k��H �����B�	��T��y�J�D#�����B ��,\96���^$�SD1[W@����|�D���n>��b��Bɠ
Z�K