library verilog;
use verilog.vl_types.all;
entity Engine_tb is
end Engine_tb;
