-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MdmeGZLyyqbZU6nx+uJBRS9uYMVx4Wun449JL3V30sr2/bYopPybXMmHwhjYK8jWbGtpQGQz140M
IZT5ONep4CrvNe0m34hKZksecfDD2HMmgF6aO543+l+SpAz+Neu6YSrQ5HE5x4LJPdRhna97Vw/r
nrXC2Q9QuRy7gZ5pj81J7GmAI53qiuKTIREbfC0nlJtcrWJJ2ypt7WiAVNGIMuG51rwlS7NAuxhq
U3xzgpllE/gtSOa6BhPSBWFQqDSiNvkOZVRChDMeDLCvUjs0PIo4ZY1i8MRZkt/uPnb5cOu1dG7T
Q9wC1JzlyCDRJC9s8AGioYcJA0nK2e5heF0c+Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
okPtI/ztuHODeW05lyTAkluIvSHYtqj43NZqG5d0r4R3+u7wIKvHkgdp1dypY6ghvi9vm4u/3wqm
gbJo/GzaIUB3HhKcfFHuLXqYethIu3cUEdhJamfVpwnECUvbQLRBGR5U6o3Pz/EYrjX4jfXuveb3
twIv/C+5IYizudQRz/WeHgoX3iR6DECQNI1xKg7wbtwkbr0/tIXNpb7ElxSSJhc1ZMIHx9dtUU0l
aYSQqmgpgomxIJauLPPjvOk/lZrNyfTCzFv0feSR4TLdwnzpAPyH5DaeSlbhsI2R4MplXn6dguQK
XO9qARnhxVbviEFMoRBLwKgVEpyt97UJTIboIoO3BP2+rcIHkZ+Gkd/E5KElPnmhNT2BEw+zji4k
ITGvk7FntI5cirf+K/a2XQsgA02VHxRSBGrkGpbnEej9QJvNYA1FFZPOL5BBNIlq9kPwUTfSDoPN
fYD3zRJSk1QD51WjluNKMDt2mi7hMNy/Vle7ZGHxiWN2EqO4+U8Jn70+vzOmDhqWQcm0fez3b7IR
i0NJTi1FxULRmNFQ5hom4efGUFBi/uLXNinZxZjCMd+0zOJvQsrF9fk/kY8Yq9oPB3Chn2Zf0rqg
Ifusy7qnU0Skcx/8+81Oq73Ckk4mBKQCmYHvxdtkcZ+lSjYIujmTVuJKNokIBpMOoVdoS6zAzg5Z
yO40GiZZrqgtEGKtCHwFyasc4IU6UAj4gXotVVQYvOy8EHs2URLY0cbQCFn3jdCtqZIdzq3nc1yk
2qy5AgammMOrlIq/3SppgU5/VRl7Wf7nFjTBNf1kW50END0nDwO2E5On7pZlIGApLwaq+UQ5+/VJ
kJDOzepWPItWLpBziFY+pLxsE0RmokXE/3Bw6KWrXLJXgtdyWKcU/K0KAoBVdmxBBWaKCihYAbe0
0X/BHrvODbDT3ZK9Am/tndQsNKsCTzcTJOj2agZE8IpeptepyKWw0YAhmlXKxsuWzFy5NiuJQTXX
fMc7eo6nOKrGH3jcAdIu92Vg7lmV5lAV5jporGWfnRzML63iv4oqEfO68vOBnq7yKS/cBtq5Jakd
TM4JTd8c5Fk+jr6hQdWudE8hbg1I/rydwp4l/Djs0xSH85WdWYymJgl6b5UxpeUkY+4lnYWQknWU
2a2yNwxWq3JJ84yW0kqZRjkwE0SU6pBcS8mV+z+GqQ9u8D9D8Gd/gAnOTIlKHQP3Gkgh9VP86nXG
VddcnlSO90BINTr0BwJImTEwZmI6zRbLubJaP+3nwYIgXkdlDdvpqIiSzLlxRYXnJAtBRE9yDL5z
3Ae4+Orw5Ytn7PImGft/is3OmU+WBS8e1WubHIzkeGEwq+gr80BjSdzLAgjKzoExtETUl9oAQQuf
ek7nWaVd+BPBvwmv0/+snSMSAIgfIsVsFbZ/SAof9jAKG2HTFJnXBexnoCYswfSQ/WRe3oUTpyWd
lc+fRW1EnzG9m5ICMqmiGdC44V1TQOTULADHj3LV3pbBFB0yzVH2cg4IU8AYd8Tk3Bj3vrW7CaM0
4l8cbQ7EkWfM/nH4B6Ox5ptO8Z8PVIw0i0987MajqrVUr2+sonFOvCDUNXSPzu2Zzke+9gnmYEBo
KqFPSCX6Gj0kg2mB9aYcWFkD2MRJ0ZL13gR1vr73Mii1vUVQmPA9hmrAnpmaOUVRks7Et2LSONlN
PS2Y1XEOVraVsJAkg6DJ1GD2eys1p+1X53zyyYelvbSx4WYDRYbnWrCsGQxzbahFsWw9vXo8jpCk
BrX0m6rzZojsOhH2tj0qhWMFec7lg2QPT+4M2+2C3tyTX1tatZN63HYEgqsoGbP2jTBr2k5afV4h
y5RQ1jiJVsXsFwhEW8BepJmlHgi134jUkGdKoLCbXGfvK4Wa1iv2ZG2JmLRAvUYriUG7QxZyyOrh
I4Cw6b6x886t3O6kkSzkn+GFUwTL4I3y4bcC0DUrBBGpu1BSYJGLjKJjos8yss+NEDDWDe19JKFn
fEIz6oVVFgQLFw0adAJYwJNwvXyfSMn0cH2C9N3N8FGcGdXzUuueVqgtXeCTj5mMJAqevpb+M7Zx
0fN2/Sv7ZOESf+Rglq2MXL87mPTwNfDshUByN+G7cLM8kWlZlhEmKx1xGu131mz7EH0ghlNtYgdo
NnewEYneiglJEHhVtgHtYIa79VYlJQUXbeoIAxPHF1q2xJUSwL+OuWV2c/jhnFFxSLgjLoI4c19p
qPEWPlvkKlz5JaoNr/MVPLrFggm/usn0M12vaI2JhAj/wmJE9N/FeX0ekX0uHmn1icnIXoGzHbR1
FHKtS5h/6laSrsCDjbg+Dn5Ul37movUnyk9z8iDhC7hvDAPSFK565lOpKJJX/9YGRaUkGAzYBgx4
2zGh2ALY/RFPJOj/8jk6ZDATKc/kHJbJbMVBYW+J/giExey80tTQ4LBcEp//fOQapQPLmK/nigd9
Y1Rb3buIKUrvbC34KLv0HPV6xD6vNZwl4nVB5fshFTwb9vInD8zmwgraIgPfFp3QgE8BX/B16Omw
3W83LPhaQrQjAPPH45tl5WZK/oPc4ZW0RywY/sawPwdA+bLbr6AiboQacbSIxRh8lPqmpy60zfgL
scpEdYyyaCAAYJcRQ8QzFyMnlfp++1zmJCKRr1B2luV3EJuZ31+a0N+qjjKIOvv/5z7ASfP1V6Wl
33ChY3w0oHeyCQOBv7xaNolCNRB7ypG/6pwB0kXJDtuSH73q2uSVBC0OddErMEFKJXb0pjBurc+H
qwClqiUJWmcNCgUDHSggoyua709GJ04ONKwRT7v/lbPYwUIw+i+wpbiOwGBFpx2JevAX7ACP/vDw
kTSkL8AwHRhLgLEisvBpCbraQCF18wskV7/7DiLnXBnZaX0c2XPvYoQ1dfZjV4DBgbHMNgoC9/ba
2e2f1upMODml046uK7WhHgmBd+N8Wap/WBURCzqYd3NBJRq6CEvO8oU4PVNwc9/ck3eME14qF7uI
Dm2xSPKhqwWiC9Z7o7zp2JpCdHQ2Rc4Zn+K4wvuPtOZT7Bv+R55NEbFSeJEy42Q2rp7xYdhHL7vh
FnDMmobR7F268JsMPH47denQjR5QzQOebZvqbahMrA40W5v2PUnLDsLN4C+uqGVWPTR3zAnO9BOj
tV2qCDk0Nlp21vGPSpFtfQxyX3ub8J2lz7d73l6ulOB3RzM+ZC5HwjGzFoDz4RMjONkZpHK7HfU5
cXQzUtMCQi4YRwV/4QVq8LOAtgJLSnBO7YM3wrVuyJTBYhmR+vUY7lBtEBCC3U/i/kyGtkVKo1uY
P0s8pPWIE4EJS4oBEDplJfFYWKOEyKz7mq7NMfyZre4OOix6hQd0oVT05sFD40AwCBEueR1oVxEA
UqfPoc7goPmsWS6O96Fgy5sSfxwSgNhLtDSyEf3m7EpZCb0JA3GDlBFykVUwA87NsE0xbsG2ptyS
zhTPisSutSQlbD78Aj9eEAVzg+5Hcsou3yngLQxjE6YBSN8C9nxFPkI7DcOGDR3/B8AgWuWFqCAV
j3LAQh/fexLwpVqQ+mvek7+bgeTc3aJciwmMSm4lWPbNL/bAnfbAtqHBRpS/4GI/suGQedpmbMvd
4Id7jggN6pRHcMbZywOmP9QIWZGMyPw3rbOgDm76HkWFJlW/3lusVcVCcc863KEphN1uV+2Ugjap
p2EJ+W8IAkV1E7Q5umxziIXYw5e7ybBfN+xQf8RF6uiToP70VJeT8afgGkgEeBtFxC8uQP/7K/KB
BESmbAiwxliHDONdcLDaftaj5V/dFDluVNFpXQ9MNi9yhwfqyzTv6jN6hprLvPd3/BAajprU1u8P
J5EpaG0nKm/xuMnjQaQOoNVJV2AXYo3jJeOxkZkWqEJf0Gi2uwbDUBpwAjGZPqxIh0erWw/yzuy0
zthOtiV74Q6WxRaYEbicK8HRZqPnRoBdc7UJLWFlTGXNxJWua4NAg9yZBmSAXaabVO11JVX5OQq2
ZUgOwlPU1CFWtkiCsOvotcSUTnUYEChP5j5xiF8m4wwC1Cxh+ML55TyrxUJrpPqIqvlsGBKYr6/a
VfXVqXITNpfQSg65iyuI+hXT2eOlHnIxRs6zOwoC77tXtT3u2nEE3lbGPimWyJjmryAZjaJe7Lye
Q3kKxED6iGXCNnU4gWHPTey3f4e8zdhl4VH/oOLQbzfC3LkvbpIgx08hfzfEDg/IYCdwuXcJtER+
qCPw2IPQPwVWmUny1W1AX9nRlqP760OWehOSm20mZFVMkXaAkkDPBGrKxpGYasYbQn9yH3oUZ2Rt
+Tpqt2Le65ZzeLvLDrR9wdPPLa/wFe+r7H8qGX0rrPTh24IyfZKQZ5C8MSsy/6TBJsocBViUW4fW
LFvN0hscBw9rm7wcw41Kz8NsVofoR6Ha0xTG5xOH6xR2dw/0hP382or+/JLN+kPIv23KkQocltTL
smkTGbBVuFM0jg+NfHGXxmPd+aGr24GpBWc4noBCr470XX1pVYir/Bpr92HMSty2cFSC6h0Z4prM
UC6eFeLfyC5bh0Ov20/DsmDl2lU/OJXO87G6yVgQrhresZqhOAgRMRAFeL9iRJXYIExR1HTB6Kw6
GRKfmtcgZ17jYUhx75T5dZYO6wz6GPpnkOooBIfOabcUKT2OcWclduU1IOGIzS60wIVQ5yqPzzlF
vc3fhQBUjL+ql84Vm93vw5O0o87FbZIeW7/YihddI4PPhc57AtBLt6A34bqlkZJE/ySDwXrFAz2e
02kbWw8R1WkasQvUqadsyEZIQzkmTbYKoEcFbMH4SJi3i6a4vR9ajUOO3OZm7iwmf21LMPyPKpYm
Lujk/577HObur7IzdYdii3fMLnJ9E+i9EV0As37gsgT0EqrWPsxqJYvhxTpoojQuN1O0oeOMmU3y
im1X+/6KhEoO7kY1Pmmyp+PqpFRDKmVzc/6qakoEtlk9UFQgscL7zi7slhGXL1XH6XAmiJxy4wzR
/31KGuL83bfEpYBm73ZAmfo3HWqJzTZMrqcObvvlJL66kpplFyTgh4GVEka3lZDvm47R+tMcB5vP
U4DnhZ+VHg+LV0D9XuWDwR3G3j8juG618m2EMAtNXzFRD2ueZnT3t3MA6axYswe0ElTBkdbJDxBV
niDpX2uT5/ayP4v7CAB497SoWlvnnzl6fwy7CXV/KiREUPmmssQ6AdvtLg0MU8hAMHfqEkAxqUlf
CQ438GSUvM40v+fXSgHEDarYaGWFRB1Aua5AwiZaJSTzk1BQnJwYCNB28c59MrBItmVO8m95X0Cr
DXCryv99dVrffgrhFCwI80eA8+bcWODl320o7vFWvApr/KUi3E9z8m/LIZ84LkvVOLU1I9gR8S2m
kNIRHUgy1HHz0BzVDs3fx4CoVAe1JaNQMRzoBDCmtipeXt3E3KkCSXD85y1QCUSecXyH0mHx5JM5
WJyRD7L9ML8zE9dk45YkbdTGDpvAWog8Lu7eA3bSSTMwU8FX67qLCWcJlvGVMLEvapp/ibd0H8RU
KCJQBbO/kA2mUh9f9S09b338Spr4onqkf6eThSO/f3O/esHJ+fRRUpna3ooSbXCGLvG+ilf1/j0P
cmH1Mzs2Lqdh1gcsrMcLRW8DN4uMaJtE0vD/DKY2gRTd5ruNDFEairq9bfltpITkVwVQ+5fl450g
DMyYYVDAiS9CZ0bpHuANTe0rzADSOyoZwwaOnGOKmIpmMP+N5gpvAPNVdA7KGEYacuuvjxUtJe9n
2euvR3jHy3DzFuYmRQ==
`protect end_protected
