��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H������N݆��Ȗ�����}������XQ�ǔȀ�wu1eH��F �O���6���5ig�a%���5�Ќ6\�f����^ŶG\{���6��5	��p��S}��jO�@m]�;�ˬzgv��4�i"�d-Ψ�C��2�g�˰i����xW�2���g�~�E<�?Up��%����
���'඼h�{��3�ThE_pסsKVJ�`�j�#{o��{OTg��T�����O2ֱ���"���f�9Q\�~�iT����H�U���{b)�LZ���&��2N���-K
|�+Q,�1�צ\.�	���lMѹ�rpV+�,��+���ױ��F%��CNQ!��艼�D��cX�&�IE�u�rˈm�;�2�B���ߏ�W-@<�X��ݜ+Vd�n�0=}xf�bfm&��]3eu���t��յB�	+��:�룠l��1p�a��Y�9�r��q+����&�TDt���/@A6Y1��LJ���{��ӫ�(\:��d40�n�sh�<^ƽ��qc\+fe&[X��Ea���#�F	Zd�bF �V�%�\_߈:��Q��v��o�L�G�pC����g�Cn�����j�*����R�͖Lw�
*��.�r�lk� v��+����Oe*����2aHHt�����9��Z��vk(�����"��/����H>��#@���n�?�Z#R�pHUzGלi�/��y�D{��m/`�VM��a(q�٪�"]����*�ޡK����di/.=#��8w�%�TO����Gs��M"�>I��0k�3�4!uy-�tUQy�9k����@(m�B`{hW�9�i�6�U4�d�g��H�o�L��J\z��'S�zmP�s���$��9���nbӲa8~��v�P'�Pb�
�d�e]���Q6j�V����ϐ����Zv�~!L{��({���L��J���Ql�6�qY�y��cQf-��$8��F�'|QM��j��%�ɲ[��1�� ���G��;�9$I�ڞᾊ���7d�lq��{Jؙ0.�N�Ԋ�堎�4ȳb�J�Kb�p�81J%)3����K�׊#��'���)K��[R��we��,�Ki�"Q#N�c����rF�����)0��=3���Ք�a�t�e�@xL:f��:��5��mP�b�<|�g��#��3��qބj9��F�|��z���a���~�t��3Q�/�zI(����D�����O�<.4
!�l���1�[?�)�r�WR��M�՘쐤�=WT���T!q��M�x�+�~<�y��&���1%L^�{� (�<C9�ʍ0r%�]O:X�g�2����l���u�7OR/�-OR9	��ݎ��+*�gMz��~5%G�Y0�@�*Q�O͕r��Lx���Zu㷽�fJ(�p�Zbh:ґ���qo+�m����Z$�'���1�V`���_����yn��-K�r�a���S��I',�e;��Ⴄ�0E�#>t��+�y���I��|�ʤ�굚��}�k�.�dX��͜�l��`�d�b���9�xu�6՚.V#W8ƒ��C+�v�)3�|%|+/�u�v�>=�'�Vv�[����A�j|�zĳ4y/��L�5��+~7�T�W"��1��ڔ[��jq�+�ݽ&�;���q
:H�$0-�G86�G�P;m�q�g- �&LXm�D����;,��Nvb�lCo,n��ش�͓v
���'��w�oVBW�TLw�ʹG*�f��-6Ƿ��)�z�|Gn��N�j�}a����2@"�U�h����U�9�)����.�)�d����AL���E�ʣ�V���V/�ǀ`oX>��r�����i��kS\�0�%���kQ5�A�ɊiHS��<���S���f�ݘ �c�g,���e�\0Ӂ1�����c�#:j���D=4BѠm�����'�(e*sbM}�"~����K"�V#)tAq�������.���h��۬s#Ko6J;�8�i������U�����K��$J��
�/K��Y&`�[)�� ��*\����G���!�����=0֜[���h���K��^�ֳ�U���H+.r��$�����jZ�N����ח���1��
�;����s��#������>�aZ<��C}w[��w��H�#+x�i�y�pw�l��(��.��
�3���\ͯ �}�k����fͧ�mƲ�I]�:���(]�hr8�L��z��;r�Q�2oS�9}&dX�Eu�۷�+��Ԧ>ѣ��9�ks��&ڋ�yI�O#/uљ��Q�:���2�N�6+i�Ƴ0���JjIVw � ����SI�$y�Ohw���ҏC����E�������z�;��u����9�A�O�/��8o6�L����TMT~(�M��3caҋyYR�bCgd�dR�S�\ u�ǧ.�]��:�u؟˓���&��_v�.wr�jD+��B2.hBc���u��]��iM'm��C�ƷHtm3~ ��|����_���A�Č�TV��;Kr$h�#9��أ���VQ��A��60G�?�qc<�x��.3��܈h�奰�����l+�̜g#W��9�#��(���<O���Ô߬��|f;�3	>%�yG�d�>�(Wɚ#��#��3�.���H���
*`>e�R\A�B���3]-0G?�aB^��m�i)��҆�l�ģ�4�F9�=�,���Jnc��R
�zS�$_Mg�3�6J<���i�6���oe(��o�t�M��hhB�_����/2�3+,o �`�V�g��s�7��h��2G��S^�d�����K/���B�����<��$e��M(����v�w~���Ae�l��c�uaL�*��zo���4'^�Of\�q��_���޹8��@�W��g���C`(f6��,0��U�V�koj�@�{�sB1��	����Y�'��i9�����- �3�?�O�
��N�Y�Ӡ�kP���G�c�@"����.}���t0Xnde���$�}�<E���Fnj����a�wb:Slj�S�B�#Oo�@gU������@�{u֯��tg�k";���r�A7����'�I���#x�[����� /�*�@�-��A�%r�^
�۲��i��nǫ��k�Hx����2��Wa1����7�%�ZD�~�
n8��zza�Z��)d2�wWP�j)q`��q5��f�ȈKl��4��7C-m�,K<�n��%�q�ed����x���sr��W���j�>�/�4
l�y���M��l{1��M_�T_��d��1iP{E����c�q ���i�^��Os���N�����	�Lf��b3�~�	���:��r���u0fU��ޚ	?>�ה�:+*�`9��r�ٍ/�xC}�)��	Y�,J�g����v^i�SN�װ�Z����x��.�Bx��=�K����<��x�� ��]��J��	���i�qG��8�N;7k�O����U�%&�X�h��z���@s�#�����>���v�Cl��~�7��(�_OB��b��C#;�,_��1��T�_(^�kH.�����S^�Ls�*��w��ԗ<�秫k�c)I��V�P�Glpp&n�݄/T�a�ġ�9�a�CiFO{d�@̑P�k	v�󽶈F������a�]�����{��OrBz��xǫӹU��$�6���r�MtC�C�f���5��W
���"�®�;����\�[9;!R"M�B��k� �.�N7���[g��t� h���LF���c�I�[ߌw��+�s�s�K �0�*�H$�w*��Т�Ȯ@�s�c����7�{�֪5�~H>X���`��<M�0ܝ�BL���a�%yt_����L�`ʓp�T�(��F.��9�b��tL��oi��� kBE�=�Y0=�%�SY����K��Lmc��m��g�&PWp�Wr~&��hg3�4�MP�Ê��T��]{G�1��R^���w�����ډ�r�`
r��#��Շ�}Yf"��5�pu"T�M�n�J�A���Z�O�g���st����Uר�;"�0"�O�E��K�Q����!!U&=��[3a��\��R��+-z��U<Bd�Oo��Nu�1$�jR��X��;3/ZϿϓ�l���^\�(?��F�ppށtő�[�����.��&:~~�M,��%oA�b��ls^@Mq:?x:��T������J[�I��oYROEnՍ~v�\^;�F��.�Ja�Mf�vF��'�ٲ��馏m&�M���2�C>���3Z�!���0g��`[yj���t���b�~\�"���27l�yA[�ۤﲫ���sg'���e�����s�4�$��뉯S���7D�8�!Û��R�'���zH>��*���I
Z������k���f�PD�r�^N�I�4uv�AVS�`'X8�AE�I/;FI�S�=�7�ekILR���W����� i�Ew3 ~/�oJ���e�����p��)]��#~q�N��Y���E��7�@)�|��s��8[)�H��!AÙ����
����fQ�DV�jI�E��٬���$?���e.�1�l��j����| iF���<����֬
�����\��I*,�.o��4}�� S���j
Y_����x�A�D6BE9�C�{�d.R��?�^�I�"�y� u5#����j�YY���ձ��ia����#���E�((C�O4��C� ���
k{'���ʺ��S�&n�����t~���������,�i��AW�s�Qmυ��G���sВGQ���&�%x^���b��)N11 bӜn���Xr��{���-�rM'�#�-4G4v����	�O��
P��Tq�>aE�d�9��1ɞ&�qϲ�K�Z��=��(�%D�����w�m����[R�/>����0�y�x;.�~����y��Db:�Wۤ������M���ܛ;Q�`�wP^JPScc`_]ݗL�����(r����#=F�L��U��K��1��mo3�ʾ{���Ts��$��e@�t	����?�:�5�ʐ��&7�[\�n�NF"FH#�M�qW�va� �v23�ߝ/���cWIW ��z��v% �*�	/���1a��rr�g�β�
;��4Pv}b�[�c���g�%fr��������;ʋ�6ͱ����k�w���k�q<!2��0l
�B�s��Q�U���#*l�'�V���l�A�n4	?WS'��6��:Gr�S��I5H�-ݘ���0����Ł d����Ʃw@U��-���c�6=��M4G���SSV�ƫ���� ���̋*ʢ����X$o�M?L��x1	����X[z��0�ذ�w'%7/z��D��*�H��
�,}�(gE.,6�q�+��d�[q�*b�kC�=f�$��ʩ�����:O�B�g��޵��rY]埫6��Õ�a��z���������T,���։���;پ��}�> �a�+������}�^'�ޮ���������#�H�;�>1t��CK��/�F�$�pv9x�t����17�!�6�Ƶ�����"ӵSd[��K΍�$d�YY�h�/����C;$��8& ��HzE��<���_"�ԡ`l�Ѱ�t���)���³F�m:kߝ�t���r��.}�z����� E��+�d~-�E�Z�&{k�͎g�Ӛ<Y�q��?����jP_��җ�^f�OM��H����H7�ESL΍dfU��oV�]�����2���<^�D�6��J`��0���59��s�y�n[���G�C��������X�a���t����^{��zW.:_�#����=��dS���+v!E�\{��=X�/�u��$]�A�+���*����%���� ,V<���1N(�U]�%�󢽬���k�k(x<��.�v�C�d�F�G�U
�p_�8�œ4fވ���3�㢔�m�|\�Ш�c���aȭ®le7aևB�X��t1��#`
�;,����V'rGI[�7S�+n�ʱR`�y>L�����Y��$WІ���׍�t�D~rE��b�N@�e*���~c�?���C�؃@]��%#}_���T7��n	^�~�	���5S�7���8I�R�LYG�)O�'��U��}��qD&K�ާ�2��G5H�:*eF��#�|E��P��Ѐ�[۪d`��G��!�ۇ�L�gy���~�*E��]��ۚ6q�s`g�J���+`�i	�.�>Cزr���Em{@�#��~0PF$���i�ml*�2.����+�P�E��Z����ݹ��ŻW;�d�^��ze�����E��