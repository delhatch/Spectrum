-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
T/T36xYRShh7G2A5zNP4dlOYX0eWKJ0slT2pd0xVmJ376bx11gZi4469iIkqs5pGpEiAdufpIg9i
211Ac9xZmzpTKE0TckhUIOGkQhy7Ddy+/I+ptOVSLHJd/jl/e6rfGS18c2qIwv0laYaTO2/wujq7
28Gp0vHusds1N8dAgH9OzsWizgMSJnjofKQcdYlFq3KZxPxZwx/IUmKKKYT3nUFU4kfWYc4/DTtQ
wZucQ0HcGboDKIUEG4e8rW5ip62qDTWWVw7NEyH6i6ctBBwD42+yY4UPe+1U8tWc6c8ZTMtnzTbB
Ow3nbb2iPy550RtEh7NPakeued0zVSbm0wiSow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24752)
`protect data_block
eXim95Sa2JKcsmWs1ZbWPUQmbwrn47UUlnD/7si1miF/O9Dj6nyEQVGwrDObm4NtDCavmgKZ5TN/
W9YXL2WsUAiJ3phWSjEGarBDMTndk9KciYRf3DyJs2GV7qu2Tu9Jd+y02XSAXpDbcAETAjQwAHtX
OTydUj2wY44DpYHwcOyxVfP/69ySirtCk99FqLaOlDr3p2Kpae0b2zRU7WBqHpC8Soyf+R1rksDC
sHkRn0w4c8sCESamGvPevPJidnsgiWJ9zS1RgErSUrDNIzVCDi6ENWJwdzG45tIRfohJEjrQbklg
W6OUTblOkpN4m9l0RlDLB69qOHVeGeXGsMh7k6x3jkZVPU6C6J8AXGWcx35JC6gMBb4R5iy5G73+
czX7u+vcCW99dGqOijgDqViTuHR2OqAr7nOvUk4n0n/cb2f3pVEP2lpjaTBbqLWJExZbchfynpxA
us0yc578kGDS3ucq/qZDiveTWSBHh2X9q3whh+auq+C6zx/6Dgbp4Rklqhp36f/z+Jadu1bjZ3ny
2xN0VUkIN6tNVuKSoeUutOHOLaCo7xf5+5/2trC2lxF0ia0lUikKS4sxePPodAAzJYTz6eLqdXb9
0QsztgpMXLPX1pIDRVc/zzpilH2sC+ITaJXJ/YkjrrAq9PQ9XDS3w8iyRm7BClRcAc9CkqgLDWZQ
U0/6D4uJIbPhrTcBNrR8HExUTfvmHFMZvBdMmZSfWl/XZHhz3lHWBESN/1n65mNoJKMb+EuZ5Wpq
9jHLD3oI0hDKe58msxvi9Rr0OAGrd8YGzPJb7FhghBsRuuILUI6xMl4XQ60jhOehO+5F/6ncNjMm
pzh+z+EleDP7HiuPaF9efJyRIiNWa5jPQ+R7K43IQwRAADFd/qvLb0SzGiqIYAijCVjC9SVNCJzx
tWC+/1aMNzfdULJ3i+sRW87tuD8toclRVpDbD/TsKqleNSiku/HCwhNIAp2jsEixUO4j/XOmN7gm
wSqqHRrm26+5AvJyCvXItcf6sUrBLj9if3r8I6tnhX0xp3gCSWZ98kYsIfD4ixejpr2TnX6vcuy/
aKYHx4EosDZHxTZ1UgKbCwQDkv2rqq0eUkPiXXTki26+/2WbyqsngMectJJWxHcyQYHIYt+Uep5j
ImubbW6Jps3oQar1U+BH1L/L3bGsAVmvpfhTN0B+7vgOUL8klCmY/igpoX4XSrRlOANdWNHiJUZw
GRU/eaX0bF1sLkbaZb/xxj8hM546vbYsTMknnoIgpYxwLx8Lexgiw+cQ2DBQUKZGLN1imIH6fLuL
oH5K2gtYh6pas90mnO9IQI+9dmbNiGqlDwdeflStGm5L4S0PxyWRvOw1+Oc5zOoVYdvcSXEs4sZn
81RMRPiQwA9gSdwpC0TnL8OwYcCaedwpwwhrotp+UgK5NDE36xgNXvDe9jJSDDC9OVYuTUixuJrc
QsRHAQ4TU3/HiWMfnKbaHg9KTqMkhYOQ1ehiD9EVwMxJTjNhS4qPtGGMRLLOQdPngS8/lfgKqkGx
qNjV048Af/br5Csa6Du4RTJu+mZdjMDn581MwcQZjriV3ZwqQJQLEDj03zCTeW3rWkJyAtK2/3gd
2PX9od2VSDyzanF0HiDxWZpahgx7VN5HV91CqDRSjdlTGJoJLDhCA7U20Etdvw4W6k5RL3cFnk4z
2I+1B2gATb5qwWT/w9raQ74pUeUX0bi5awFDMTaXm1YdfKCvB3sD09jSUgv0gNdryjtzy4vfx3yK
xcoOzFfdT3QlNH3Yi80EGxG4PMjuz2ijVLKiQQxQVQNY2vpQylYNNQWXXO6g/Cll0g7zDXgHzwLR
MaEivfp22rNGFDspKxllByZMUBA9LzYl0hVkP9uwR+mBmqyJXBlUgOEYBLsjlpqF7Mm6zUW+6oR8
TU2rqBoDgsx8XRbjOu7AkDl8iY7tePBt8JZ7giVel8SfB5OZr+9DYknci0+kaheqvNBUfa4g3XgJ
AH8adWhWgr/6oPV/zJ4Lrk4Fm2gAJSzTyB3is7mzE/ojQy/OIl0LAuc/T+pf83dVIBJicqjh62I4
oI6o0u9vOi8G3uRRex8EV5uc7e8Wz0MLK2Q+/X3ZBMs02iQYj4W0pDpZYFeJ5EH4C57XEfAq4BSi
cQpgGgpwO4jYQHkLypF/Bp94mlu7r+fdnKaKpLmmvMB4ePl/qDK/4I+7hi+jTNcX60p4iTff0mxX
O3Lvtz9FDO/DzetpwbOvzF0EbR1u63/GuU748x0O55dr32lDdqGLxrLMbbCOOwEC2iHwXJ/YNrpd
JItPkPvNhx7LDUiVZ5XOC0gYzMw3tw0jExMfZwiuDP9BUmHnHM2DJm/aeh5F012bbRYEftmovNFU
oJmDr8TzX0ZFQo5Jh0+1JSkPW/qpJurgmtdntQruPim9o95gGVyLlYa65yHozcIxtGoZZLnPoXzG
cHjM+X1O17Q7Jn2Fb9FaKQu54FrUjf7llLp5rqEUcBxQGHx2nV5oI6nKH9GnzttnSdIoDJpWO+ZH
oPX0Cwhneas+uD1wF91ePcqw/DnmWyFpol/5RwPJOHpytAurWSQQdG0eMkaASu2zff5+cZShuDuI
PtOsq+fWio7UAYc6QTTEFme3ynP6bJXluNvOssJ15+1Yqx1yPH0HjVAgpWeN8a+o2M22wx9mPkNv
yuT4KlskQCEjvFTa1Utk4nFlUWFpNYwy+PJop/OIyQOcpBO/8wmRusn9kCrzh9Ds5QQuBbCTmId7
MudEdWaoUNQ1tebgWM4S1vPN78Dw9JxwasT94Ko/H6Gz5vZ9STcTYazM2rAkNQPa5bXqIIscHX3I
dZ7wvm39k/+4PvQ0i9dAL5GsV/liDKoOBkM3BJ33EpYYXzq9Qz/VjI4HLmHu3LAE8O8b2ElXnFkw
2JyRoiOTTmiS49tcgXEbvxff2PzkXAGdBNVfbrW4Jow6WDHjrq/N9geJumslRVfu0rRMGFnmRZWR
XFOc9S+216Gu3WAM8jLM253cBbtqjd5J32v2U9wgI3rN3wSq2SLUvtxQwLAlneAW6YPBL0WITEF4
qCAz1Qa41A9tPabQ37ULU3R9BHSjx9qUlR+1RozCrfUit/qAWQ9NnK6RdC3USOrfWx2+vzoaWl9x
Umv3E6XhXs1D6I+OtlAokyuFFlzIPqvcILSAdLdW/OTvxrv4XuZjeqZsnZ1tKmBUNO4ADpCpH1rE
G3NPSqmG+6u+Yp6bxPxn+kNHdY+skzXMy3q6Y6Kt/LHYOBEbJ3Ts8FAm2BNLqcNFGShj/hcl3Rp1
y3FSNPrApXqs5THlkmwvmLhrOAyP3Eger3+dUQ3/69ll027/X4fNYbgygU8BaRuLchjChdn37++s
TpWHLjgZZFMWPcgWwDsyCW+n03ZszwUy3n95EQ+DIcaX8yLeoKcIfbMvkP7mX2ApElfWY8/fiPP8
MF2Hs1TNbiXeaYTyg1S+J17rMxc7BiTe40PoKwbeiLVW+nPar3EGhQN1zkcWhPb/14quiB8hmT9k
PzA1zts+j78WsRB9fNChcoGja4pLhsSnmkAnChAAZE9xvhl5GEbhoxC9G+0/FgHkY5Q2EsmVttB6
DbEZPguaDWvuDvDw77d3UtrtaZrPjKiRVzfeCzTai7xPtcfLaibEK1s4n4lY05lZvF2PtxQEOSHw
OCqNidqYZ5V3f6SvD0ea4RU8M/0CIMOTbUvctLnOuTR8h8jEhW53ilJy37iqADR3auhKScMFrIc7
ZbmE2WBn5PU9Dpvr28IIGcX+feGmvFVzxlHLRXq51kDH0dcX+XTu9uKC/y5xdp7cpg+tGMUDr7m6
eiy1bxhQbGWfXDc0aVGXAmeWT3rkC+rcsSfvFXR2qSudGFwScTdeBNzoKsazxRd08xcZlToN7f/a
w8GazQ3eMtyee5/yRVm+S/hc1LGEI9l5ByzBRqmWqWOupTdDz9LuFcSaQT0Xv8QET+rul62qxUhq
EOwGfXPUwa0PHpCXuGbxKQLInjH5WYvNK9vNEOHVE4kv8xFWIGFKe/Vv7ehLYWKnJYnYPgURFCcg
GQYLdAjb7WwA4K6+mX5Aspc8x18EAE/tUu66Bn5iTNRE4jsiumJj593o6nENzaD5nO+KszH8LsqZ
BmR8/GzyS0vfMU66VkJdU3sWt8CjWnSc59234bra5Rr/8SFXKiaN7543aqTpXVBkDviYo4EJgno8
ajX2tjPMg2LdZ3nb033ue5Q8Yrc/ToNZn1J9brKtwM+AgRQXi9ioReDsQE0V5siC68oE9aD/Lm/d
HRmLZK++RHpDRsToMLfRRP8+OrXMpam8DQkTw5glkmh810OQ2hd6ix0Ntgg4Vlyu7oiVkmraQJEw
dlntH4XZo/fBkw3pZDiv9LLWAFAxRP7A5iOqKp3s+QzcxDvqE9CLqZzYFxQ/C2rt/wh5EV6Tp1Qo
PIqxTG3/5OHlz0M9//FJ5HomCgngqU7D+Vp4dALtGo3QXVLNansDN/yCDCvjyAuWQ9BK6phFjmZp
D748mq4evmE+veTML7Ws8gD8yCNLIT9/saQQdZ4cjkdlB2EAYg1KV/hjzRY/4RZoyzB2JwOrTEDG
p+VSC5F+58KCu9pLP5Ydf31ONFcRCBSoKOYIOIb2V13fosOTKYp0lg1bjah0FHsztsbNiPlAcN+t
WOLYraj0xUC8tqdiQ2mor67zZKXS09FodbLy43kaS6Wu+z37P5/FBaO0nhKZUbwcFwREBkkF4R8r
Kycj2V/uAWh4/9JOJdgLF9PjcsmErOyQVHC5gqkgiAeBAXzIOaBJVDKnvikr6+58ekG33MfKzKu8
oQWJbOj8rThwlxbmAkJvttjW2qblOxKIGOtj+hnEEvQ9gQFpyfMOcf1yPTQ9vAG7LrhN3YWn9SKK
X/skxK/sbif2S5OMocBwz+RPGrBHtUyXYL2aJZYJAHUXJFv5SfD9HVL5yH2JPpXsmyOk5j1eDUOV
I28mR7ta2ornucSzK+SmP5Thdl0opqQnxRF5qxTGiccA8p1VIJOo7q4CGTWoL+27NzKHLM5XpAg1
ZI+Mxq89naQ+IYee7p/CPOiBGXgghWG+lCh4V+NUhmNJe1Ob2/S7j1nydAIeEDn5yE/G79ySHyzd
oj/tVbYglTdV4Df4rnsD9I/wTp5Ji49wVLFDmnNdqB+e2GqYNPx/yvJRymezUVZ0e08Trs1l5S12
L06iWe2k1wc+hTN1Tan+Aurqy0zvQsdZy1hhn55BnAklRgR9udVQjep8TFqnYh5sx3IVQ1W+1tvq
6keKksOSNMccXgOKMhjPPvhoWODcVO9K/wImuLyunkKpdb9aikdH0Gb+Eo6zF+hhKXhI25Hi9pgf
KZyAcGmTE/Qgp1dyScCIWvRR5P/1OmQZqEOQ9QPsi9W78n1WwwzQU7pUI1uVZOfIoF/aK5zpDyL0
D9yxtpqTBR0EwhCO30qSqQ3SJRvtXqLtCMuBFV2mVMcIXJKPX9m28FrfBkn6Q2mTaSzZSLDfInQi
ow8cz5bElonFvCMYTLrWS8mMamJK5jOj9A2sL5gZMWylvB385eyb1ZfYJm+3xWTdG2YO0clcfdgC
Z1c17Do6Hoc606rs2PNIFBtGc8Is3Z8Z+/MDJjt4qso9nHrGfyN0cGkb3rCIHVo05rHIqZV++vKu
EENQKDSGtaX+QDIaCJlyLu+LChFzzqfi3R7J8YVckqyeTrGSz8wxeILFx6X17ntboXSt7UsOcMhn
EvVU29UsL5NVm/nXE2gLTw5F2ourSRt1DvHQDTttROo28HhzM4KLsdn4cJtUK4c34efGdomOgDUV
1Y1twj57BnIIj5nxeXs+PV1YODgtDyM2iVbu5Zt97eoPm97lqmFXHVGNbN1c7ZY2VJYUrm383O7q
tcC/L5updp+OL1uKUvF/HVzb77/rVaYUKO5aPKbv5rBcEvxmcm4lrEc/kg87N50opP1auJKiUrXH
bmz8DMWT4E8dJQBKRNEy5EBWNuxCUFR/PCuV18kHuKR4g99WAGTd1lNAhCgotD6GxWRSMnKIVDd9
DPV9uaaOOrQ3FWrtNmScFd61ki2TB5XUjxW5xpUB19zmbQpJydesXWTqRoMxhInncL8wvs+uxVK+
L98FzvIXpMmn4+9KwvUHH6DEapKExUlz0yIIUsUJCSEI7HiLimqvIvgOAwzv5gBgk2iKkSVxDvbz
JqQMR1bdeBMsMpdIBti0WkrAPb8F2cAMp3/ytpEncn837X/9VruvY2rbLki1vfCC9OZughT7LWZR
Ku7mjj/Flv4PSBwgDJGKf5E25DttfIr0M6mF9FEhrRiqIA9CFBg6QsWVEYBrqW7wl83pp94XcZlr
wxbG2Wx48wMSFIOzLaSAZyT6ezUqJd1stIf0sWIhI72SxV11NBvCDmBxiJjKpXBh+kWgfmUpnGvb
Pyr/cgMzCZiHbAmnedveN8NgLcVkDVjQveEuMqs7XJ3WpIUHXka2djdN3oaFCcf77W/ei9P+1mYp
m/aO+fP/AfVSfwSUi50uySDwL/wMBt2/i5Qg3WI0IeWICMkOs1tnce7Pq2QT7tO/MyyHMCmyPtID
+AI9c3Od2nQ84nc4MBpyKST136XQvsgSEtAlVjyUHFC5RcyNdF4GNxY64HCV59c9Zhd9V3eDZTd3
uSCjk/va32Gt+jDMHsdBGpJiqCIvewASZ0NXMoR7tvTmQ/jRNJtpSEDu1CGTbQg3EcWgOm8MV2In
F59alh2uI6Ed2Rg3+bjUYyCjLzAU2yGJW7bpWY9TCPQhr+QHJo28qnHdITDUt4XekiNzLDCC/9CE
hcH5Ph/7bCRrzNOqmlsfQ5ozpX983XBKO3R3no9I+L1f8/statgE83ix4kJ2NkmW3dz0levlfiSk
6g5VKGjeCYr82p8dWZhkzjpfVqPCUAF/2UzIZvzh7B0oTTt43qM6rbJHfl2BEgS+tRHmGGGPj8Hk
P1njVnLcDPn04sAXkKD5F+2ryesJVQOkk9IlNran6gt2jr7XPEo3F/ISAlQPTjXUXaO8ViVW70z7
lAB1oHATs7OPf+BqrhpOoGd+NXrqXVF9HgvqDpoCB4CvTOzjObddUZ2VWdcMCOZtB9V1WXEE/lS0
rFOyfrnbEXiwaaSpRTTtuDRZFPDBc+d5hRmAqnSurQTNSnQboRLB3kBd16qfbNAqH2v2lIHbJQEF
YFLAicsctzNJnDUgRm/+JYgK4VLvRQYFfR2B6kdIsmaJNLtCURgwdH9FxWwG+OzH7hXTL6XFykFJ
hpciEAEkwccHAVIiHyaFEa40zQ35w8E3noUFGPBQbFB0+kHzf0qTXgypyGlXOQ6moeycd19QHN19
fC/H3Q35G8VrecLZwcsmxU83UKJDBedYg0t/qUpr7jZMkJ7zStjTFwB+KIsCzVNtJ5BVm/Wnap2/
rl/KJH9PImKGjEsEEPjXcHr0nYO2q5rTpqvp41ErDGUJltta+mkZtm3HgTHXizpOHw0Wua0031ZF
IkDkp42AY0jzKon71dsI6k4R/cAYR1MO/dggJ8BTnCsxrgNL/5BaftcSH6VuONZDyBHqzrONUxKJ
66FuJnj0SR5X1m87hWdU4jMPKAmZX+ydawpVR/LxzM0tlyELvcYILernycaMDCMPOJGbODzasW80
m0NBHEasBA4y+mDU1h/QILheC9ZZm/9vlDCr96p70jlLLb+99q2KgqkMPBzejOG+9QtI3hlAJRN3
PqrfFqbBW45q3deLW/lUecdKIkE3AieOGKSe3tUKG787aBs3FPJjgRXB9pYIxDaOtGw1KceaUYuW
YWCUeq8MCKfdywCBTWvm1mao3pzHI27RxPq/02Ggp/dzFw1f25ga5Pe8ClrTJwh+6IZfgRz4Iz6V
NOQlJaPo83bkdfP5EqapKCsRabv/vjKlPvcM/vj3La1QbxrbZDie745KI0eLrct6hOsj1PwH+az0
Dr3NURaxPQlz4HNLa+nIBIyq04KPpqVIB+BfQQSua6RpsEREsCFWC48qduQY/fbJT+38as1/aaBE
qIyqA3bCN7h5etPHsquXSzsy5uMLago8Tb/0Ckt5Z2ePdQNklK18qAzC4oLHjfIeK2BOZCU+LHI/
CzNhlub6Im8Yhrnn2Qln17CfYbzNEzIqBEd/LQONVoZuf7AmBFXC/OSZI2qx+gjR1TZxKXmV95Ci
SDXPvtRb17C6rbkzZzAd3Oh4qCl8w2Cip7dJPOt1wOrOgIuXkquxfBsC1fdinc+zYSSI/CXs0alX
GeG27rzGmGIugGaVIne3FBV+orsxd3XOvrSAuYuY7wf2Wuzlpmw+TiykREbZiIw642elx5cOwXpp
38Wz76op3Kzi0I71yKL5mKooZbFgBNnDDAXVVHZS223d4wVt4hF5R77dgnyp1zrquLMpueM7KVaM
qv9S9d59sREsTHQMseQo4/8GQj/rbPHcqkm/YPFv0uD36IYrvv5/mRn3t7jqxfsikMDb/oiemQ5m
paJ9AMOlALaabVc25Utzvd9Ll+9KEgd+c1Qet4S9W6ewnJGoRtD8w/nyePkMEi0SXH/rCg2emLbX
X08av+WVB8seuiMRKj3PDT8/ETe+uFJj5CByf/pqSG7e1ZWEEl6iq07tdOjEClF9YaMOJE67M4jL
4qbgD0AqseL69h7sZU32fGhYCkOsHoPrPAT0z47jtgu/BKj7zM6FLZtpi3tXkozmCokX/k02EpMK
gYWQIEKNfgcVocRBXzsbIrmqtiQG2u+Vf7x+pplvd1dA0grwBDxL2AUWLYXfpCVqC6OFDC9NxU0H
x39CKwFSYX024m3Aay+14coYA5o2+yItthOt0NvVguzIB9YZIK+I08Hl2Yf/nv0o02ncb32gmQaH
nnVMf8sG+q2aNNZE6VdZ6xs+r5IVultjv9lMKa92hn6kO/Vphat5ogufbeqcWnd3h9k6+1AJkgp7
v10IF7zFH5/Vd38uWsN6QQePOv2BLhbixgrHnt0hS+NDqCOK26mKSTKiP7VfBm5k2u66yFXfh9FG
go2ktKRZqfNSRb6xFRovuvN0uz+P3YEz/DUDMF4keR4jl1Eg1Iy0kT4YlizVf9VDr5i6F1jD7XqL
dmjp0FMaq98rA/WzsZrjNPw6pDQQ45j+63FgMHeAyOQ+jVNyKHmK5824D/vQCJhGz0Rd87Yoe/xS
cu/higiQ/c31A/DC5oWwL/lbWJ+9IxWDfhP8P4x40keweMZlUQ3Y1nqRjy2SWc0/vYTSUR7kLOf3
ijf7iFVxPB87OJ867Uxu2Mq/WjIJc8Z9tb6KjxeJQgLC7NFqGpcOYbnFLRoQNjXzf467tQb7z0+V
dhxn30lW41FfgXS382QQjxeUq1yUJrezOHy+YDS0c1Jx1c45Ut6Iobk8OlVLom4/E9Hucv/YyWJo
HgUGfMfMlvB8KexxrJ84SrS4RWFpRkb+ZQRIQMKqQFbIqH6sC/5g7aJ+Mpa3YLTp2LbX6/Vma1IG
ctdx652i0GqiXrrWFwGYLbX29mMs9SmVwYdUpsOKHBWVoFwbq7Z+ykcmgNC64sj4Oa/a3A9/jF/A
UKSdXnMY0tCeKeXrgpkOS7HpWQkM8LEq+3yE0JBq5o1umxDHMV4lAV+nCh+/1t0toaHC4PY/VvHe
QvD4/F4ewZ1ScrZCQGS+gH6TZlr/vJzQ78mZaZz08jCV5HcjDibMtCy43CJfAzzvCn9s5770SNAg
u2xAiaTqGG6mhJNauco0Y2xiImS7q8dc6rBiirspv93DAEW6cvdeHwbuRdy66qwi2y6KG4dv1Vv9
SygnlaRhlT609NaRTQl4hFVdB7HtmjcTZql04TXZJO+UOeILlTVhSJc/FWub24LvJDLuLgFeoDO3
5Yx2Wr0Sc3+DvbHLkl0uMkYw4ddt++JtrhhdB18peqmQ1VCvuzSteoleBezEhkSjyh3tf9Ufc2Ms
iyk+eVvBh5C/sfAyYeBkdawSUXlZ0PPQeGf5kvgoiVyks9neohgEVvLKdt9c+/ePx9R1Pyu+Hr7Y
3xBAADTmjb8k8ObBNbf6XYlGLM9ejqyZuVy2TmEyebCnDzwFNipppyUvuOOvz5czAULtxXe/09um
xDpExtfuagMeI/uBPx4ccgDTGMIPwizgs6meUBU7rOxZZtDjPjd7YHPIKCLpD0rhCbhhWaI95IBv
Dvb6cWW+ie7onlgP7YdXKA+C6tW2+dTam7IcWFDtwqI5wMLoqbNVcOgbFKBtwrs+kJ6Bzn55o5Ay
pHzEiFceNH2ewlSeg9Cw299APCFLOKSNw6+isygGdVTGtDhNbSSQKMFXxomr3/+C+PkyWyiqlati
9KlVFZ4T3z2+D2mTTaN3A32eV9UoNh7tOjAb+iSQkBu3Y936QT3eXYQkaBsPuEKhQGAi0IvpRJe9
HV3NxsJ7fZMIIxRI5tjuBx0qiQ548QOjeMYNbdEuIPKeVaO8q8JsdZdRg8+qyxNnrofD3kpVOXyI
Z+QJ8cq4ofDIkhevF4AduF6DPD72bc/KGzZcrAHDsImyq2W+LIZM6hYe2VPpmHpjgJA9lYR4SLe4
PG5bpveQRDohH/HTF+r4nTtSm+pRG9uSwSNvJxHizUZroeadj8r4OtHFzEiyy5Ti3BCW8NDxh/DM
sE1ZFY2C8mLmF1iv+/Lt7cxQrDsL9H/DT6TzoJ+o13a5A2iPG7FeZvciUFT4+XpY2F8f/cJ0+Qu0
NMtPZf7d0Cg81DZKBPqKJIFRV0Q4jmObW3RpTDAFzupyus1x0KchDNrKoafHETzhTNfwykJkgHJt
qYcULRMswerE5WrWncJZanouh4wVVLHPotvMBVFnqYNYH/wG9qHhKOKvXOgz90lub4GbH2g8ZyjN
jwhnYqSRPJHt+WM6kbrooWb30GfAte6RxqRXONcg8+ehogo0A4pYR7wQ2LH+9XiuOHZvfNHdpdqB
g06SS74g7bT7BXU+0Xo2wkF492zEk+6jVy0rGbHNJcBRqYN0yPX3Yjlr6LMv4Xkrf69xcyG9htvM
lfB6t7Zi9O73O+czLWK2ABWaindUbuoGL9EilR3vq+wZREQ55S6FdY61XjdwJ6FUpu6nS6k9Eiqf
uPnYDsMgbfOGx+bGJ6CPGu+UdXwc956CVJn6BPqaiAyx8GGMqu5m2EvYjjlDz0mXJOK5bpmk/fmT
uKqptPz7vgsW2DBAhor/1g0AQEJcn8Qiv4vn1SMdwOtR2FQkSz/P8JoQWxYXa2bFKZTjyJHZTy7W
bP6CttA5KQjTzbGaFzO3DRUew+1jtTDNcYIDfWPyBp5tvZe2/AUoMw6W26UTpV1vYPb3PdoRHdtZ
QIQgT8Tgh/8iPIJBK2gTLVnjL78pmH5gO6ZvtTFRptqtMFSNZisuvBGS46+X8WuLISVZFEvkvWnJ
M1X6oMIBbT/VJfBYbumnaScaP1LbGOs41ZZ7NVKQKuaCxWZXL7c4J/Xkf7V/xlG/5l8nMUbCMkom
nBDdBZDvMKHHijtECUmsRmuK4tGVgmLV6mD9rKtogSRJPeKhR3KKO62Nfz6w3Mjxf2y5QZVgrqpn
S5cJ3SKCNM8DkAUh25YRAjs4o7hiW4g1kANZQL+uJc7HKjVF4jPELA5OyfZ6VvkbJgOozquVJC2t
pN9Te0kze5pD3YdSXKuVNqjwIkih/6rpW2ahdNZqrCZ3rGHbNpeJ3hvaAVrUO6R4fwtDAcZQfW6T
YO91YC8rdT4VkdkZH3sRNC+j4aJmRbx0V2nCuQbP9x88iX7F0e25XygiSkrfLiD5KhRyDXFSZIUh
58L//1e/cfvh3ke1vid+qPdhSljfte7B6onquUBScbkF8S/qSBi2Jy8HlpLro4NQqSz1nUEM1bn8
6e25CCnuOiQRGgTI2FHIvzYdOP/DFh7BiHbqjEPdyvG8mjl2gAmgAWrVqC7boS2ZPLotpCuIuB+n
1EKDZ7yrw69zXnucMA5UFt8U5x6eoVQfYLldth1P1BdRrOU4CcoObLBO9vMahAeSVud88bEN1ffH
gyesYO0taLfmGYfddbO8GUasqsU52rZ2TjHTxbflsu3dLN2hqjkDtRe4HAPsV18nDBpp29N+Feru
dFtqbN/Tx9IhzGzuiwcs80FRJSmSS8n+1HLJcfvwXoFeb5of0yZAR4a019Zvk6K6r0tQnlYkbRss
coM9u0SKrabeH8akPQXwOD3x6FmZ2elGMEuxgQt9p111ewDT2H0fzDctW3VsqJZ6SV59YvqCrO+C
iG5dLBG96QuWBiIdOIwq55Wemxf4CrLENh6iYulSKRNZwxGSJeExfO46zPJjs1bHtLzyGo8rr72C
VTzW9DzS1WIKNytRfRJDwa8fEzBv5PTjk/PCfVBhemQ4HO1VALjX80vW/IEXjwNGZLx+kTZ31k8r
elc+DQ/BQudzAsurI1uhVocjHm70+bPoFEDRszLuUOL8Bait7joOFLPlfwx+lBBzKzGAVt2SpMpP
L7SYGwxmf4jHxITFgJvWadOECxUpTDY2R4wBxeafNpNJa7cztlCb36oGwyzi6Z1qEHzeU+XfRLZF
rePRZFXB4kiFrJ+sgkzJyfIj5b9pY11/cNQcKSeP0YOcLJMPi9qwgY2c3TKxe25LcEJ4uZawvkRI
32gs4zwuB/PgHlnMX7UAvLgyj8aG0qXTV9rOEGq7jxoJlLO4I5I6zcT/gY/4BwpBz1rTOtm2ljXp
YVX0PYv5tO8ADCU202PxOPpl5EpQFG51MjZ4XITSnNoOHxUUbIQoiWhyWweN8UaPhCUqdxgvQEbE
jcF5otHxlMZrltgNeiMD30yL0x+Sp6GRpz+jMXjverImWMSft1DdJCpUmpQCYz2tJflJAeNIZkeb
MPFRroJbTAxzzCmF6IxgG9az2seZ5ZLOoJax9IznUygub3IBiF/S8FSGKcz+ZrRva77kOGxVMgU/
wPyRblZkX7bPFKCPS5KkRrSHGO7TUkEHFRbx+3PvXuCiXbN9cPWTULvgk5Q1wvoBszjhBDg/WP5L
+rOrUTosmZv4TFkr7X7PRhnj3c4jd2ziZn+sLpKtx1RxnRMjoMT3wMoBtqCSKmQ+gQK6QWecOyQH
hXBfvD/MU1DvWr4MkjjPKOF5Lin8nsPVrEvPzA8v8qxTuJJvHQyxCRedvJQc8qN+k7KfB6HnVbNA
0woKyvtA63R4ENyHRANXDC/22+G1YeoflSRHRVzbAnw/msOhUNXyZW+nIJMNJEGMRrAEbCRHMcpw
limxPZTKF2XjIYIWFEHe9RwIgAqjYT3ukeGn6LS4oswbS1yxIdRyGmVgaOu8aVOba4BpDsmzlumn
PsWfM+2xuD1lSRQD0EFny5MxnagHsZdhAv90uYHlXtYMc/jabOQvmFEmDH5H1Bt6mUJtVnnpFKMR
usDNRq5SS7i9TZZClQ1qCk7phFADOfflvyA0fjXcDooceWiJnbAr5rV+TAwGRqOqX6zaj1TKai+C
87+cnJ0zBBX5AQCGiYuJaXwXO/JXvo/d26rEebTqdzHo+4xxgphLKXdb4fwhlhlkA0eD5Joz5gb2
4mcIILk3AjxIl1rfvgzlkNxZu0Ha+0dT/BZXVOQdbToTsxj8e6s4abQkUzVnC1/p3fdZp65LS9+A
Q9HtCdVLU5icDoltbu0rsSWx1n+EUg73MLv/4mVXNj7CHI4AY4Je+j53K6M3ei3ybO7Vdx++Rwzr
l5v+PJJVkgKsn+1wNo6uM+vryM8mVSx5a1MUoE8qri8A/iJ8lp7BGBeGR43JaPUH1ZLGK9nNKJ5W
5EXfLR2gdLK+h3S0WgxG59/Lsh6ve261MboMg8K6eDb/YBh18qWoSIoHVK0jQxaxnSLNUVoXqfvh
AyC1hpIcgzR/pO5H9dXlo/8+3iSVEcjgaVQ1KdO6c7xt01iOk9by8p+5q8VnYHKcj1iZVoh5uIIM
gKX8v38lnxc85W6yShXO2wZDP3Hg+YcxOCrKSBB2JlX9kGKMn5V630CI97AW1ZD6heXuOOLRXIoC
2nrFPLRlE9EwTyjNxS05OJVO7NBK4EGP8/CCKQCJa8JCkiS9ZjIKII4sokpPP2YZ6JBN6GpWsXiC
jCuWQ4W22ZBW3+lMQ+6XNVf9/gJg+jMEbkOjo1Rduy13Kf9SFiYShKgzZHrMqZeEqpX7g9ZQ+K0J
voIqDYBAg68ViN8j81ZF8WoANsEecVcldO6Bk5x3Zls/rGQv45E/+vt6Ub6mMsikBOBSECkvRAO+
86Vy66P9MEw9ieiQKWduarC0Dvn1b2J5i5q3/jq0VwZlGtGlKBW5S5TOZfRjhReM4c8sH+QAEFp6
qP0g+PPrKGqSLLUU9XPQtirwHb5foJxEbmVi3MklmJFQS+wgP8oI7QJwtO/88+IeQG56jHWlX/Fv
mugOX6cSvICvib7M4LkPCTlQCpdgqmz5/0xYX1EmRW/3AWVyutphoNN5vYvkwKwe8Qe7a/dVFMP9
/TOIz5PmhD/j7DfQoaZqWp+qR45sRsOV2w1AehjyPY1JtRJbumCA/dItcVpk6X+vVYPOajYqTyRh
nc5/LoCaW5vagORwN0ZLfwd2OUGees7WR2wuaCtXHLBhSDLmxjpBbv2XB5i40RWKg1pYtCetlIow
io8CnQHvleYvSjcIe3TKsi9UttUNyKRwVqjvQThYYt+o6riiU5KZMMjYRLLAgfDMFabbF0saHZUH
4Qhw5TDfHOUBR44QkQfczJ9Z6ajhwKBd7MSZK2ItgB+rI307e+JcyBCosmg0rlcbSofbkQJfdIBU
0RH56O+P1icXohVKcME2Cx3jBqoNt0L/zrTexgfNIxWUeF+12ATNadHX3ZaF0bPgysWmVoqgxs4B
YrAPmWDJTU1wtaIaLnlrDd+L+YDguBriWmUXEmR74aahBFh8c0xGi5MBcfXH2uie4h8yRolp8//V
kHovWcvWxzGxItas8xRtpN3cMXnO5HSh4COzoqEsXYRX0nqQ6vWcW+hhYriIXjZy6fPG5rdoa0Pa
0X/BuWRVctyfSIsgR6oC/rzaKPLcf741FA6Jzt+96GDCsknsgCX9ARx281RZ9MxmlmuiFjTduYrI
nJf96DYiuzfQM9S71KSq6RfP7kcBWwhbRm3LMfdi8IXfm3Nzfui34ZoZFDqcT6ONPaxSiF14NkZ9
iEP5u1B4LE7b7zEValBjmcF7jD4CxKb+geB3dvZ88I7/B0BB/LyTzGLuwGkWDcORfePO/z11yTRg
Z2MWKx4XDQ8wRb/gMGAQeGirHpXvYk7Aq5lSrfRSgssLAjQRGD2VCVP5UagfZfoFkJaKnoiIvfh8
FIi5l7efCCHkacNYKShT1QYoafwBRD4O3EtdGCgZURnrINWZHd4LckNTStOctURH/FedXA2qo7UB
oj8K5TsWZdCZGfCuIjDK3oZhucTWHpeLM1fbM+pLy8rnp6d+uDfnEre5VGOZyMbWptzgeqn6L7B4
Hh/2cdIvisj9sHZkeq9wjnP0mVBDOqwjVBFqRYbCgtKdrOmSeDTPAsGu6GtmJN8YkbiAZTfLt54r
4lqTKRD0FAfWwM8KI6q+dUvm1YKbHII8KWQSnnaW88m4cWgp1gK0hb/+TTTjrzbvimt1xlsjvg7W
sc0OwhUDn7Bc9MAsmRVpApKdSBlK/rDjrYZUT2CXQiE0STD8sRJNmoSWIpSVnSycQgzC87ZFyQtJ
5Zy+nVtLAXmBSbiDxCyGEe0ibf9AhrK5gfqXpGGbiyDlDavAhzU38pslDH9FhNrfQo82vJBdHzwp
t35dT9aTjzXEdAtBo80Ri1G26ZXIQSysyNv4odduhEZpbRdwqM2X/o1hgZmPcEhxvw1gy/xElCa/
Uj1JKP+nfPenNlepEQBitZJ+CWefbplrrmWWy85Fx6i6f8qR5mYkhl38VLLkjIWf268OfMnCDloF
9VGaAYk6X+8+7QUiPy83peWGaU2tPUaEhnhDHpArxQCrNjEsFwHu6aCDFQUfGsmEjQJ6HGlPGp8N
yatIVw1UFZAcmXb80I7V/4sI85+V0A9uHdzxZlLC1HeYbT9jkop/67wTdjpg4tAWfprM9WiUckEz
m5mEkIBo57uzM39gVo3iDrrdbK2DeUdW0i8565M483q8nAs4f5+om8lhBZfoE50c3KZNR9s35cBU
cwwh07hiFQXCYyDKJ7KRVksTFr4olCas+FAwoVDZVuwguL9QNyZ+6Ub5d+E5nE0+X7+2rFCwrjFx
9w7sYRDDwTmk+70b2oT4PmERpoABcm5YwYfw04LAnXIROcmiqd7rpzeBj7YkInii7MXA9wq7/HeI
CpLp46DM0tI3I7eVDIS5DTKC+J+tYGydRzmKqBCWJRcnFiLUOO6A9LjrRpfm/Qy9CZZY9CFL92cI
exX+hD4os84/xJFdb+Bj+oX/rW4WFkVT543zxIBQHLm18rem8Ylm89MbiguNgcvcTOqUQrykddKo
oz/wJJ0fh2zIGQASiZIT+N9AIAo+Qfo6txIGnMfyuX9OM5mpHqrvFEQT/qMkrLohKn0eecSSr9Vm
Uq6Al8iDBq870a547nMC7NsI8kdsR4LEgzgXdAnJZYXtp+27I3DAgRWJ6ychKNtIVXNr0ehGikC7
xXiQiJVjmP2NN7n9hgT9kMC4e2TqAcg9AqQpFifvS5fOnsQn7MD54xRrq7ZpnW2wwlqqaZrotoEN
w1BgN3w7OGtRcOLnfkra2/8FwnHGn87D6OXjGYra+GVlt6OyLOdgQsrCB7l09gqavFJ8f2ggSaTU
kNFBAwGA1WYesCVBe5J3Txa389bB0rbzbXMASqkneZHuvB5F/ZoFkcr7geJ5amDmcFc+H7+Y2Rdo
wWnbMbHcNLWqCnntXyfSKzIS2GHon6ENjSQO7R3H4gxUwJdMu95sYoZJNJ6S622d47rGrBk/2VMB
uO36a/LBXkTgRNqjbpoNs2el/BuMwqIuLTBJPDlg+ICJwRoXnIS5bC5kWruwZc7GwtwfwsqlrgPR
Czdq+1Ji0JLdZ3FlTnatph6RBs3pueJfCyi72KF6l8M1sR/iTKf0aOqjr7PUH+jqNSJ5882MfJm6
Z5Lsno4e4vP8G3j0ppK4VgJ9SbJgqKn9K6AnmgPnrbAgFigP/+2K5+IbNfHLl2ImSDP+b+/+KxWg
3Fp9tRyDQClyr4x1hYcu/m7Qc/+i4vBOVBMfBW1A0bQ/R/0gfNG0EofZ6PqjnUqc4d+J3i5PheL9
hnRyKsdNBJinaBUA5tHEvQaGTg6EFm6xiNXIlK4TCCCsJNjmG/eZu2xXr7CHFFpYJ2osKXmAVZsp
ppuHTjx7JDONaiYCHi0NogZFElRAjmKC+iRqhBt1lC6XKP8mA9JHWcGD0F4zNq3f+x1vZxHsYIbp
9M4rwfyui18KCckktRS73yjkGXqm5oe+4VuObFiWkkxbEW+xl1EUEF+ZskSFDWR8mQ71TYMG4NU8
SoMgWyG/idKQISmBRBMwbxpyhtHZJ3KxyWcYcdhNbTEux5BV/JNvjEu9yFyDflHziJCPTzdZFOVj
ws5p3GJtD05KJE34R6tIFYcyEqIDEbcRnjf1J+/ytWGs8CYDSxrYikYZ4Nf4r3kuvTX9oq6utQpa
I+ovenTrKIg7P0ViGRpxXIhAh311z2lC3APIYKKoe70o65ckXoFW5j1tH0ELkq4KrMJmd4lFEB9P
tMAzht55bo1RXTBD1jnXZbw1rjelmBkVdz69pdXa9pNuczKBBfpU+HzzjPe4hSsr/BLPj4cqro8u
E3/VWI6c7K96ZKpRy5dMTW+iNCbgadOVpyKVCDmZVl0uChz45FHYFgkCtEtw9JnQgw2Amn1G6Yqn
k+CFxIaDfz3uN0SeMAhnqb8K1q3wNT5woF5EomtAsd73TqmQMphQZ13RalAn2lk65Bj3597NdjS6
UnnchgFShtaY08DWF3ziu1iGu7i/TBPI2W5W/5EdiUcPAIqsYQRL2Gk6tMurx4auRsIgoJIy51hX
mJfmOBUtLnX8LnUCFcN2kOwoHsOoQsoaQBShDBA81EIkV8yHcdI6mnN6SBfFFAR1pLyivbRj7oER
/AX6HeoQrud1MMg2kW8vhmoVZP+5J5p7GffM2E2xOoDSC+xnvJUw55+368uHCjlA9bHMrd0plFgP
75EgcIsgMXEedrrbRfiMajOc345lNhtWCCEmlg9qsB1c/A5JE0esou3+usEsVBGIAm3rCipfpVDO
DY4bAFZN70TtIFrUxVaM1gBNi5FsLvImh7ib25ZHNyPaQivr4GJ1TRtVP4sS0+TCYl7ZBucw6/cB
664YPowiQIQuRyAnFYBu/n3hPbkJROap4mE+SsCN09meYZOBvDU4ylaOER2eSWUF1EcMVMo7vbdn
jCixzPseEoNvovTp0pDlnxB6BEYwvUKADuB/EnqgFbLEewpK5hI7P3FSGMvI6nMrIZG21ew7rT8R
ydV4gLdspunT/FKyeHIisVY9DVkjjhLOc5Gbs0mg39fkPWE+7OUpZfEOdsciXv/1OfiJZg5Vr0H4
5MDGGxIbwaf3gmGspVg5uKtINUQ8Ry5lD+XDqmoycR4wqQLVfyHOK/oE1x332QZDvkQAiJkkNW0K
qgJ0EsktRPwT4BfTrgjKGukjLeNdwtitHcBQ0x6y/zAHfpJJdIvtwD0BXdxT0ljX3n97MyTSqtQV
cXP42uiwang2g39iB4Vq3tkRsEilswIqiGFHDGvmgLP0az6Xet0P6TryS39kOT/Yd3zYCE99T65u
CwZJoctyXEOROJFt9gfprnKIlDEzFlljJ0lnbr2ODqIF2FP8QXlHwec6v6V+jTrKFeaW0qJOSjOx
0d6zG7Vo9PyX3hSvDbX2AGTTv2sc2CCMkvGZlVzfpIGKiRThfErcFGogt/CYj9Tyc36OoAuXfET5
yQmewwCUp8NGyLcXY6iEx3ZARACRG69pC/0wY091hYYGULPfgX0mUpPv5Ak83wcA2bU+SNLMWHAr
rUJqcYQHrtJle04xM7saoYS3OqiSkceNjw4j6YZx1Q1ywwWMb4N59HGRCwui0jKMOpwaTnwp0etV
+1uBF1dNSz49PpAJUuoI3xtepBB5NwvLmK8QKhTZOcjI74WFsUobzMIKpEY+wlE/huH054pl5yNS
pkiOEjGoreqt6R0e2fpiKS2lJkpsZRKjfn/lMFH0lMyVL/mGBxysfSawHrJ4wi+sT3QBZHOHAXfZ
yDHa4MpUC2YkEpz4dcgCpgGYST5TGxggADSjgEdByNNtoOp7fU+yyV5fLYT/7xJ1WzPa4rCIhI3c
j4yBtGRMCPL0Cd+rCypGEZBlqs7w1gFDZhM7vKcQW+DAcZigZGVtjIFEeyfo0NLVCKV1dKeB7Fzm
Xpl5VkKTOtkv6ZnEhTrnSu6WAJplvyRghKmYtIAPg95L1biYyfOfk9iKENE8iorE5Sx8hTzP01kQ
GGPHlPz1dSZbZGcfmeIhLJP6nOVX3x2wOhjrgwDlpzmkT1maEhqD8O//rBfEQ+gFPf9uoIQ67pXS
jmvBmkHNXEhsP58E3NlyWWIVScpjcjvIASe+6s8NHK4Pj35I87jqrp2fd3EZZ86X40nYhknr5QYb
17DpqWJyhGWvsaNLPNkdMF6wtjiHw2Tj9o+QbzSq/s6mSRKaGS72ZGlf0fWBsyK13i8GgwetFfJh
RI79o5zLXwe7fNHMOAq9nhRZlX07THp+Hfa179sBxdQFnXqRTodfXZr/sWrZ+0EL8GbsUwv16O4w
gOrUGpRFDeKKJTvLIB0S7b0Yy1Z84T2Wab61S/2QzqGNqgPOhCBo4YaI4enAD3lh74aqO85ETfu6
jAs4ty1SAoNdEzkPm/NFbnJ0dUOvNfS8CZb8BNPlV0XNzk+i0jrqHURsKzf2MlJkdxf7qa6mJAHV
mKAiflZO3d2RzY2xc7gt2s9YqXYDTHt5Y45wvKkyia50tvIxYvH8FCr3xMsjVBTiFXEOPjLiAP1L
0NpoozutOxcWzjr40aUQl5YJSvVzsYyQgAy7hctFwI4442lnML4GGOXW1WhdEQrvocjcdOyjOSwJ
3CwZIh/Wi7aTL0kArOefLSDcAl8kW/fiK7OSPmdRfCwpyzh0ksVD61jxzxxlUubAcbsOsTTR0f6A
QAXnrXv4hb2yY/AWw+8OtzREPIApUlEsaa2VjM1IZrbg4oZ6YHUMb6LKp1U7bq452mFQ9uTpnDVM
t3K0PPJsLEIkp987Yq9A5OgugPDXUDoj13m/hdIxgqEK8VuVTAllP15nt1xE4ZPutRzAMg6F6nTE
DVQl66G8DB73VMbIIQmSOANMJxYgKGoOHy4y7ObslaVyZyHOy+Gsu/48S/4LDpCnA/CP250oZEN/
/SOiTlhJH7jC8IDf7Q+iIIHHRA56qggHF1SoaLQnWd3zacuMbLO4Gb0xJfm20u9XJU+3oS83dI6R
fqJrY7E0CmOm0SK5gSj3eGVIP1sUuAaAHFKseKJG81AZmm059301C1deEZalpJytg3ZCwkbQa6YQ
kfCeSlzm9EkdqTOUgLKdC9A3thPTFKYfHhNfM+E08nesznX/mQJLXxleN8AbpqyPjm5u/9JGBxn/
iqQVuHFf5y5dENnirUCX5ORfNiLfyqDM6gygXvRMJD5Dfp/4aINjtKXCVlZr5m9VJT2D8ovrDGi5
LXmKwHko4aB4zU7H3G0mqYoVqyYjLsbuPZrxiJlp9chqelf0hx2f/4xU5h1G8TQ5IW5t/VDXixT7
v8Oj6s+pUPYFnTQgg7w+Ln+8804h2cnYbjgcX0L8sjJn/4C1yEuv9LVPUqCDgFf0V6lL2uKALIvy
5m7skLhoxDAviFhGRQIWR0kyXU5JCYsTsQ1jwu4GC18ns12EFmVv8vEYnzLKt30lWo5jSns+eW4G
wNw7WYZLQ9erLn2xdfvzplbXCZYqBpnBUfd+BGQouJd5kCkSU+6PYdCSgHcKvt+MIB+Xj92Btsl3
Kdd0fpj+3CSXbgANRdto4XSwW0Xt2GnBBQsqxNOafBXTHHKWo2nVklA+BUROvLGNIHtnwjhYqJ0c
xTtTuCsXQQP5odHWL8M5ZqRL30eoN4Os8CKGAuEx458TrxaLsJn7pOF5mLwNqgBkkeHRZNsoYBA8
jgpzA4XZyIVGY3wV9ffZpXpDYs4trYCAR0sZ9DEF4qV0PleWgVQWLOuMdCCIJAKwvXmgUWaB1n6y
j5YMhG43y7q0F4NikbmF5/m0xxi8DSrVc8MJe9kj55kvqokEupW4Xh2Beqiobm21W4xRVMWc3Ie6
teGMMiAW+fX2pCYwWTOfqNyo3WeW4T7rMk5j3Z2JuY4bOzxmfKBbQA2/69wi+Ex4cEQq6xzeNhcS
aQ9VxBAphbeWuoKY/ymo+OL6rcjBBXw+ifYPZxfsWORVgkoZJqNbtj7vhfkkDLA4akLUhG2JRMVy
MPGYid2CI1NuHrJU2Ye8OV3gQQekKcCuKvFLx8XZtCIOwCsnC83seF9FrI3QAwm5r510MFF6r0WY
clbb5g7iwzQyW+QvG3fKpqgdhlP4Q/GYjopjDwfJEuEnhDnyCtNr8JyCywnu54LWqJks7/mN+MpT
MoLVAw0rOBzq52W2fbSb34SMdJJZYeIozSRc1YtRmvOHiowHu1Ay3CW/ILeTL3sWcyim+b37psC0
LVC6WIjnhiyPcMJk516RUbEI68DbFQIVtwfBP83YZMSlKoBMt/39DST0RZA1IOdbU9UOibAfjtDX
OwwBDQZTF0FsqWFkk99hI1Ln2U1GuR3BgRnb4+otPxe9j3ZWOZPpKszNExIf/XNCMl6GsVEiQuTX
JbGyX/0WWw0Q3UAHpAbZQ0amkjhhj9G3sUZI14tCsKDZA8TiP7AwYk2O5bHWYPOF2A2JPXL334kr
pY3WYEzr2c2BUzHZXCiB7K6CP6izMMcIVhTf5DYFWxecBfMZOAbpWiwf0vYBnN3mSaxtmLVJZNdX
mqTMdwgOCSMqPocDYwFaAPh2Hl6c5hC9EPXfEe44f7CNQlBLy9e5YtqDcBHEAchuRQ3vJV7Dscjl
p34PWKvzxpfT42kwffpTRfm7+mbHii18Lxh8PCifG1x1XPNlkMsu1zMIMQLmb6GKedQ6pZ4+Fr+g
XwuMscw9Ygo+juQ51Qxw+Fj1qMS7rr9QktaDhVyejKEdrcue4V7xppvFfLQIWYpiHFoa9C31AeDu
2D6yq4mssy+7QMGycF66elzMbnFRhcu7UyzIrZQsnuFpH8MQFuilYJaXrs/C4mbNsK4kIabo/OpA
VrC/Qjx8NivPwxa2sKhprTYMtV844+tccMIKtBCUj1WbfWzY2XwVsc1nVHASMpMa8eV5cGW18iog
aufI/Vq6+u9OFNehPlfR3wlJPR7WrOvWGi76uqBGauRdlqJ7JF87ZVDG7Sbp2dAOmyjbk8LOY7ZQ
xjyf+JWO5sQ/jk9LwK6ssm9BpFsz4W7JBpMgLD5Rq30ZK2hltZXc3devoBktAdHHV0XZ31PvFDYq
Yofcw9qExkYQj2PVfs5J6u5tF/w8szqj4aoYHvUdPBz0lQ5rRirWKdhaFZn06UcsF4zD/5O8+6Ab
AANxcIIdsc5HPhLibghvL1bOfP1cwZQpcsmcqoIsbmduU8RlJ3S/IuRCCifGJCgl65X0PA2u+wzh
uRyhqY/okJA5iHsU6lJjhereUeg7XKx6j5grrvd0gj2I+sGRdYUZRc5azRWPU4jLvIs/munlFS1x
eT2MiC9hLcFOFtpIZwqMtQGh+b9EtWggxRg9m/s0M8xWdPsMr4qhu740sYKI+UVRpcBZxTE2soGZ
c4zVYsUGhVtaeDuljeWSqFZRN3ERil7uOBjKmg2NsfeYu13m0j/lF4ovrNr1/VIx5QMlu/osnmNZ
pjyGOE4gQDptoQYsKeCV3sY+HCfsizYfH2EBXXts+1+9g3WfvvOxLJfeiOBCE7dq81VWy8pQHJEZ
2jrYW5MIdK5Li6kzSIvA2j3erqeNh4P6zva+Wc0dBSZh3kqF5VGkRnk8bS+VEdaXrimSRsZR01HY
TUyQKVg1jpYkFD6FXftalBY8w5WeNZD0ojnS/YPkfv2VrqcHkKB9w8sNNwqiJsnCCzvTAQgwya6e
vC5w4n3T4g5uF1HDFmj2RSoSOX3+3s4J4TJHzetP9Q/dRLUadhjlNODduXMA/CbPRtuPxtpIzZ1r
6f/MU7znNiNaBERwzcuDo2yOc1G1Z9P82vnDtHYIQrJYilXkyHyBefUPOEQVkF6YX/46gC253QBw
4ZiFtXsRPjpBgBDjnxiRM6w+Sr0bBb9QZKrMm/39zqJk8y9TktOjIzJ9m6B0ezAy4O/+TbomcUfw
U86oxq9Ryih+6WcdHpHSD+ZpiiCXqaK5OCk3GAErpCzMnafe8HKD6zKzwuYCb6u3SIEsf4AS2mOH
ox1XTuayUZAwiZBnMwY/q6hbiE7t+1HQHjJCetdvqxgjd7XhE+8uN8EWCAE6Sw7RUZQ1I+7gADOH
ixodwCmQ5Dm4n34UNDkn1/a5VkCihDjsj7WdevScWuwwvFBpRSM9YT2HabdS/lugC0JUzTjm46Be
EYtE33FKuq06W1xe1/lGjWkbifFelpXpDQi6UzAx6xohi20g9XC14JzBuu8tGUSmdyyHxSEIP3uK
1VXWZ83cixetmELqOPb4FgabdX37zx/JNJKPoqJiANmj/axOrkCVBXV2NeUE215/tM9YMJVK0YD9
SbThoZ/PXeMLW9e8TQuJIuTkZm7E+yOcAZL6RDUBnEFe7hUPMDZkYJuY9hqGd2ozeuoZ9oLv5EBw
SixqDk+kL9fYNN68uOUoaXRRfBOXmPUxVGbZt47KZWayLUBtfPqB3LUMEsyMRgNmrD14SmLSMjPj
E/Nuv/D20KstEf6z4nqFyKQe+pH9bTXBawkbT74WbvEzbZzfyfW6MOqk9ZFaE38WHtoU+Y+a5DJB
diV5+xXS4eBtcxHeftsqQBdv9pttIh5TBUPwBneb2g/iJLYgoXZgY/K9Zu1RxnhzqlAH0vsGj0JX
no5Dp/BYBhIO9uDcKsL8lGUzNYt80VGV9XMHTlkzbWTW1w37dEEYIRi/aNhN9olMh3kGCq4/BI6v
54X0gcjlcuBgZlJyU1V5ODxnupr+tvsCM1AhdJwNMt47r+Oef8CORHPg40nnzHDMb08SwSS9oQHK
f4C/LqgT8/eqhB+2S92REoIpa3N3jgHDloaZk8f8qhrucRMrHh2qrq2lyyTP0n16D2g3Bha+y8nv
7deguW+Op5UNQ7J/Oa/+2z4uDbODKRiXAid3gIx63h+Jz6e8yRrYGhk9/kLnQQ4Jlgq8+Kukb33i
0o4ZS3uqSJFh1iAdM9mEI+wNRKyECvNQkmQt6HiJ7Avz1unbzBKo1bJuaqlqan5REbc+rE4HTg+4
Jln38y+WAhXxu55Hayz1O4E6oy4kpJQFX8Nh8KM6s6GqM8wfqME6GnJv3ykFePC7dsJ4p+y4RGoh
uKoCkBDMWxNu6+iGng4xjwTyf1amQoBZm/IMJajD135ZleWX/fLdy7TyNVmx6t3k1nhd4bSdUs3W
lRFygAl8+DcQvDL0rLbRddIx/1N3RbZdM5WYp8RDJIlUYAgaPZu/k0TNrmwqUNojZH7qkZC3X0nx
L6Y9F/etxBuRb8PN6PRagnxHZDxP4y87x0NjNLzQb/pZlEEPsfQh3f4ixwp9vS+E2Be34GkVImDy
+uYfvVPRmrV6Zj3rqX0oYdeK0dM2lvc5b77/7vQvLISvrYeFG5vVlEx9cYjIRkp0N1s8IMeeR4Yc
+ZfwL7aCO2wF3OYVFoDCyCTfDXNuGPFCkWmceo3PXMuLg07vvJBTOUJGfsuRJQS6Ba6byozvv2Ok
Pp1oCOCp8ZsHkFHSfdmy/MVxq6xE2L3cSkqvBJUFssZ44V8pJ79kiIX9pqoDEnS3tpcU8/5+GLx3
paQUKMbllrsHisb8qrv0t3yeqAgOJHRegq5YExW70hGJeBtiJBQ5c2qbusEOJw6Eogk4XaQ1Y4sK
91JmCFc0JEviFvT4Irmwj47gQy1x/Yiw4oAd45eJVaZ7tYQJwfWIO3hOyK7fdYCPK3U68nm6E9uc
tpjIzmaOee/bfSUkDb9Q34VTuIhzZjNjDTH+SaD5IdJv+70edLQwGRMEIFHAGTUAK1/b7LzHOI54
E57BGRuSTgCFjkDSOcfRf42D4oOtfm/TLqqFgPmsUCUd6WvJgGhs6lyA3LjaX0yDdynPelh5t2A7
8ETjuyycemjbiXI/nS/9c6deVQw4Dvim5PKwocMainKmf2jkRAzEjyalmivTrQVDzFPeZkZZ3D6U
LH24u/u/bufBSa9tf1hE5cSKNx2TPhZlFLnzymlcQiVbqqK4ZkPp5xawZscGS+HTJ1WOMEtAerWL
6NpYQeS0OcoUFWsMSi7I9aJ8Zod+JLEpTFR40fU5wX47vE3ZHK9GME7DIW+WsqAGrH//A2F07qFI
Bt5EFIw7LyC3i0lSFbfPIyRgOJUkHCE9PbD5JG+mhTt6jn1y9YfVmOwnqvOQ7di0itFYihr5/1vg
m0nkt78zPJIQohCZ5YMLaaTK2sKjRjG1fLfeeCTo1shf0Vuy+7b+AYMoX5K8u1q+P2HZ4uF+KYUp
emWddw3hTS15Kp6xWGgDKtacUC9R76ao8PWBUaPEDNtUaskQk8PzOglgovHztYyYiabZCcMKCoZs
Phi9hAsug1cNlLEID1/bptIt3HO/JFBTFwyN+p5xwAIerTCVXL4JFp+Pre5Ti4lAwLVTbuaKg/qY
aNbNHwlHkqD24nbyKU60+ZYXkzG1xD57vhWdgWtP/basVfRmv7CuWCsAP1AHdZAUiKzuCkpJ+vRX
vF4vVUq4VB52+ZKo01iCqLGjI0hio9zymYA1rhLA738lylSHe1Xe8TkMD1N5iL0jvOoHPbAh8cyy
p88t2bmDeuJuUIrXZ58v7JxumzXzt4e2VuLfcXHjkTV4Bu4//vZmMN0xCiLLl6Hbd6YR0D6wugjV
GAEuleIINh9bprwrmgU4DRNoV6CjECkxOxuPPCeoaFtnuh5wipiAUqMz815/AovkdzkoxnWGiQ5d
3oou++JnG6r2Bqet161tE1ZiulruYX+gR/SoDbNReyXhXbX8md400eYPMTcZo/yPThBJfrjM3fRz
Pjl7uFj4H+rz2tT3FoyZEAJ4gJRHnqskuGvTsoxqayGDMRevfHC6rcDX2oKo2W0w7iBXj+vpqvzG
rIl8t7bDm4R2lCKM9Sv5bS2VGRkX7RPmkMy5t2kZsx7GmHNcgawDEhZRaoblhzOHKDGAjmoy7yTv
eX4eWVrJR0WpYuNwymhfyzzPjlN7j9kubBilSCrHUgNDSbUxYsVxZh2W2n/pkuh7dovmLqoQcZH4
WFHxGKtJdGIJC4Mn6PzgSM3/3ByPZE0Mb8E6MKUsDqlBib/w9wWYO1FhQpJ7ONiq5lf4Dkjwp3/Q
2cAZX1dw/GLlmRZl1iWjHsbdDHrZBRHRcwUHcXO+Nnrm97Q0kZOWBszOUhQjJ1pWmt3D6DX/sLzs
jJ0zfb26khaTlMN3jeLJmLQwmuGWEkg9Kf5fbHMjQPM4h4GQuFv1stiaJjnk12lsRMveMI9Iguyg
aYVdVgWCVNiboJBqd9OY0BdV03OtFFvBqwaNvHFgQX1YASjSTVLY/ayCOERnHfxnKpY7gcc91sQy
JzHQpTOoXA53hUwZfRY6cld+HLYryL7yTl6f6ObURMU4Vw+VTZFVsqLv7+APAjyfADd/hDpKElak
AsL+uch0AUNhvP4xFr2HtDfC6kuJVOHh/rtW/Y71dqQM4M4Jy6NUmaN2w5OyT+e5eDidvf0+APOJ
TVcKdFxocHR2xuG8d5WPhliyEgBr5J+SpXhBuorEnSy4C4jAZTe/xOHRvJORG2H97TNAlOh/HU/s
6dtP6QDTPptKuX3tj5F/SXiy3dC7No9UZCVdFIzh6RYNDnGffONX6fkO1e//i3ez/WgjkW3+bWCf
QNvvPkMVpzrM715v45aCGtu0L0F4GM0YxGuOXqU5VOf+f9Fi4z+YTZFBs8ooRl0uBCPuKnMThkQo
2/bCIwgmdtRaxel1lYw2mwJQw/vhYDPGOnfDO+EPhTLa5Xfvk+DQj5496sdmVs3q1uT9xThg3yM1
ubYnEVaHcZ96HCt+tLhj1gKidyV2GRRskTfkMzjC+1pXeuikJepEtvuJ3x26OHOv4cuLWiKtmLNF
xlUIQvAD++DgS2fObeXx9WHLQkwijWN0K7ILhuEl8KIpP8J9wmjZ78I2Vhm68Hqyiij3fdYIKyKI
Gfh5IkSMNU/zlmiHmMYLM5WHy9C485AKGUXVVkVcFaiqvxND27F85REjSH0oR2uiKkjf6z8Bu8eb
d1K2gB7uFPGpbCu70gjl9nnKt/5+l67X3pvS6LPf7l45v/7wHAkVOB95+siQFkI7NmUDGaw7e+ct
ErBBe0rO1j9R70CrIBlcpe18jzlZeChwFj7otrlykp31Wz9/FhQ9v6K97hLB25rg2I2VqLH1RfAM
t6O9cKNnFbWlqTIVgzH9kr9kBg+VN8gdZCrq7HW2xtmyqjaqaaYjBgeYdAWK/4fT9OOeXOJGlAiQ
rOnWT/pZpVE/BiQ7QSkSFUNKbSr17XtiMI5AvDFAKlDwQsttQ0PvcoF9uOpP5fExvG4VVLrQYmv+
2lxdJZINRV2KmAR3plGaKtjFaV8IfiizQRRGE6wcIBBIXbumGewaDuLXmE2nsahs6zUwRgEmhCdU
hq3Y9WYGBDD3gBXjvK+GmXnJAJHl4FyNKMZH/hiueacD4mNiOyG9+1nu9X67Mby/GXJUwCiynKj4
mdaBaFle7PP0skEcwI6NOTsLJgKmt79kxdtBbou0s42j2UCqcIMxYatYa/z9D5RBX/BjyeQVlehA
ByZRyIDiBfnakCFHU/gQDSig5T18ii6Kv0EHSeOLxUqHqV0y536iip3YQcrRcm7bQP9SBueDy4GH
0CZnfkpjibRFm/BAqmEoy1wqm8ncB5Jw9qOUAEl1wUm5sLeAKxtRIt28pyEmpIm6xQjk2dveA0Um
KEOy+FWZ4QmwGMPPIShfoddXtCreGhn21TzdAE4I6sH/l73d4dyLHhmpGFU8bSlf7jF7iYhUIG0r
KeXiQI4G0RL8OHeu9gnXazxdJVASued/xcjbvfRUHqP0ROAZPrBbDKhTbL7m1MTl5VXy7dBPBnpQ
2x6jHqH6b8jSsa+vxyGDOnvhgHr00H177WD/PrIlgW8TwH8dBsPY5ttrBRfQ8QOUZGjanmdXRJkM
ekorclbRD232UbigXBBuFIA8IKR62/L1mvN2ihDkmSur442iGDHA8Aogq1M+91GM+QqPle/8cxPd
8cdEat7EBFXxS/j08czt9nEtdd0eqaH7ijfP2XpoBoyQyQzdJo87td1BZ9ZFRhd/EmTUKdJ71k/Z
5IjVsuhveU+MKu9PpdOj8SOFO3f7z3AaYtDLIVISoRfk5EYlP6leXn9uhX8V6KomrpU2OCwpGlQS
8ubgAtVK37hPAgHWLs4/vgcmnC6sDvTlDd0wxQTmFUYYkJMmnIzfwqzC6qXvr93C/VhOpbMOqaWq
XEqxu2bddAz2rYZfALuMsQS48e/C3mACNbhsA+4mcgj+YR8Y3Ivr6HISy9cIA0Z9IR552Ryu1X/M
WsywIs/qofaNLgJv1qtfvfOVd/q1NOb+pSZNVqWeDzXWsngyDDcIwApaZwAzh9YJ0qwv2NJnSBW+
BHTCsYJB0gIiL1dF1QI4ClB1cMAfwf7i6Qym2nFYt2B3iu/O/l7xmriyTkFlWTrLJHwKozh1DiP6
OxwNn2Yq/U0z6pKSQ5/z7RmeRIEA/Uc21HV7Sm0GyzD+FR5MqE0u8mws3dy/F0XmEdnBwZw9w9mH
easl8gdSaAT2XGw/2wV8aPlo2JEcyUuriS0aqHy7ppU7CDc3kSYmtlI6GlrDJRGaaAuWAbEJwhzx
sDkak2uj3kTwOH7d1HtLrAdRNCK6EgD/GY/amPot+Jx/cDid4BuX4SmtlxjWKKj7xwag95gPp+mp
4PbzaCkJ4HHXWhjJqVUVBjlNJKMgT+rWUfQUYOR4/EgUhWppk9WG4Ly/mF7QNcyfPy+v1za4lXS/
04uZ/K8SFOsxdjdLKoUdLG8uiThngK9t/6cSDNh9Yh/UQGXKi0Q7LlO6TpKDaOaxhb1no1VFi38P
3lBtc2VgeE0MzaebinlUfKLymN1VRSO+zVHlApuptg/KCEFKF2NPTj0jEZ5CHKUJQsSyJVNYZlye
HmS9DKSTnuv67rpVYJ9C/JVImyOgUoEI1t8rixnJpzbzu1NGQurMsyWCng3U+QV7QTnQywTbQKP8
eERPV/SgF3XzQs9VrL3iduM4j7ioDqxCdv7Yko83cK2DqbKX3/8AEaNAPxTEyDKiegA6uGCSZZbM
B7DrSGiTKXLkjBSQKbuhRkiScb6n9cu+GnwNtge3M6vx0cJ9IpUPUnZZgxbMwt2cnsZmBJy6I3qM
0uSQ5wlgi9gYwTaUY5nbdrRkECHC6btlZGl4mKjH06subjjrX9orjlG3pgkZNAkxCS1jINFrQRg1
AfG+iwttwzkQx8DNhjT5xnTWHGJIwdI1NJl+jm6+RYpALa0vYhC4YDZLpVzwVRwz0MyzTMydtTGm
lWBo5lNjh79IiWhKGJygQD6zCPJqrF9C4qeDsqV9VAdKHfnauVDMtQz0q3HJ1aMK0/kXPAt4uB/C
VGzBstcOh/vR2b4VYHmttAr7fuEjEV06gJcEVu6qK3sIAAaOnHnFdc4xrrh1ShtkUP0lqAhwx50p
INdynWxkuE70638ZleUlu8DnXAZsRoH2yAi4gXq79ptebLm44QgGiiVoXnwZw8vD2jebSRDgGfEn
L6TUTR/10zdYRjaixtQEB77l4MV46iHGgewu2lBk+uHTtnRJ8LE71nR2sP73/ORIb6vQn+uwmlaL
oZkEzpOZeCnrDI4pBopESvZ/vE1Le5NgkDZIfMuzNTVeXctbgR1J6sV4cUngHYdA7e+55ZlWlo1q
dYh6yHiFm+ngn3jfU9n9M/++CxaGJRufGPlueXVoJiotXlcSAgoMHhTjKhVTwCS8V2Qy3QlfXdn/
CbNTBGIDkUox/4aW6ygFUci/8g3w2oxK0rvzWNE+EhH3Q3IHXK+RtlE924BkvO6U4GXrS/PoI0tg
yY059meLkJypTNEDXnwlI6w/eNU4Ay6sMVjlbOe5czad2TnXCKtWCf9y4FEN4/KNM6DQ+yPup5Qf
bSEyKFKUlkN4UTJblE3LHiFSIfsmuq4jmukYwHFTnjTvXbA9Jf9rje9mpG9dn42bUqHjGlvbumO0
ZuHCBV3BidTR/syRETNRs743jc3ufy4PxKqX9paUThXrNht/BLr2jY9j2mREzeJ601Z9lUE2GyiJ
7Q5USECOxHEzRxxSg9xdiy9zNcX78lEm2yeM5XzB35ez/jdK754xbIzTwjgUT+KHFzWSjNhooqoS
J/02BvtP/2Z0QVStefNsaRirVhFhFsXVDuVpY7oBKneZH5rIsslYEvRFz7p9uc4hVGKIrQzT5qGG
DR6H4f61P0Q0MUaJ7abCLvmvX29fm64q6NG0I7uBa3jOsbk+gD81skdJu4TzOIuurXG+ddPnxt/m
lOQMBE9fSkk+DUDUG4a9ze7p07Sbtl4HS6DQpp3DrpX1ehi4IBQEARki2x7whnhEBRUb/EyckxP3
L1T11twOpCqS0Sy+P4UKgHgfWdYEqj6xoFoKnHxkY/3xgKSbB+S11fNHMRsj8ElK0lUtSzStraTA
d0zzYv6KlHcuCZRj3Q6UhckPHPqrOfTyhvHaTqPEsmC44IRPtOH9gYaGOgOSmvX47yNaHWxJ0JGR
c7t9Vdv9AEc+j1Fj5548397LpIHyphNIWfg4l8ZgWPso9jiKyIyNJYVwOCcfsBxRRrZdgUpmSzSw
yDgW8i5Z/s69+tK1BXO07Fau+H/U4P5ZIpzvIGkCaaZpv7AYhsbZlaqfZwsWGv8mDWGVASb4b6rf
GtMAn6xSqvpzF3+vvwp3yMhtm0ChSYf9AKTsUEznn1Rj5EXlL+6qVbQfrOxE7XUtYH2xRTMrVknZ
cAaPZevwsaEwAFJU45gXEM8fM1HY2VoLtLtPsmN8QL4H1Wc7t/o5XkoIM12sG9yEuYGICoqNCgNx
tbrYEYHyh9Phj8x2fRNOwbWX3UShEt2EPr+1tNZLzZ7Zw2UNr/jUPip8PS390Ew6j6Uc8cat/2LP
Mb9i/0dQn66y5IstLiai2a/fzOC30MF/1aFSZx04MwhpzyxJjj43CF6bvdZ3FFl7FpOl6KJ3ztkA
viPFatOaOxef+uzRgO4iPXRQZFhAJHF2VT7Ms4gNr19hRfYok9olC/4Xy/WUtJ3mXIcFIE2Sr2b4
PzmiHUQ4n+6tO+kexByASnX97XUKMtz784DAb9h57KBabc0Vbk14LBxiSyIUHHud3atsi7Jk3tub
I9CNPZLoyRj0IWSou0A1/q61xvq622Z4XrkMh/Ij+murb6g7ZbFA+lCSYyjUqhlXxjvj4+fb29h6
Ntq9XBGnW7exxGXF6eewgDy7NrfcKMd7D/BPPSm42A1oD0ibzALzpXCCzrCaumLjL5I4ECFguo0z
+N8lxmFns5GpGc/I/yI++jXkAitlL9gdEhpctsadIaZKFmpySC4pUoZUU1uJIf4tskLgk00rhj5G
hfEUOuw6XrJZm3a+FFTuAJ1SUjD6xvBLG8W8s8fZOLoX5uKtV0XitOy5e1cngD+ghZwyVbKcn6tr
VxuV6GZUyatD1hRcXvpp5IgPiYtuoWh6Q2iggfjN4m7KrWy4n5uDPEVMrqlVETZNym0MgVFBe37l
g9KKojyMvMYro+LtK/ff1UAt4VNrFQe28hW3d6ZbINlIxdyVYrg7e5KfFypxQVnSy/BZ7yUHarqQ
ARYxetgQCUKqNM7+t3r8thS//gQ2FWl9JUpolxCcUiwH0ptAyXicQbGxgerbwt5YrNBSsMpcZH9R
qwkqm9maJVLfCCiW/bI23UOgWzXSzxnJ9uRgXeKW6AbfXG646WWQGYGE+fC8pz65C91lL9PKDTRQ
KsCbERByfaVHAoX51kkQ66zzl0mE36+gipoQ+Ii+PcCqQ/axRE7dwL/S5s5Vu2Snsx1wspNpWShJ
Dl4Uk9XLgP9uU3INWtPBYTk301/EszmWgXtkcGmqimUJ5sID9eqbTP7DqshjVM8U6xYvREFZkvZZ
k8ZMuomIGCO7d/qabC3UF1H6mFCrnlQZzHGyF3RJu4+NOlXwvF0jsNPDg0YfM4itakgAT6rDe9nm
3JFlV2YTX5ksw4J4/TY6X7HIH2qAwR7bM1FZnfX0KklbdyBfwkQHHINji6HUY7wu0JNTpYYAORuA
Ctzur48lHwws+9QtxqpyRVuEBYU73rhmKOU/uvWuohkAR/OFqT0DOsGkgTxshrkgrms8mX3PpcPe
MBqKJAudUz3JYr8GAtdxaM9a/UVVezCY/3O9CfB5dv9GbLQ+fE/PRRbhcYD6wXHBTxe6XkIni41e
qsUdTq+hzj9/ZabOKJuCeTEe4U4LswQm38uAJ9GttediWXdJy6JUGknS4ZrnGjzBwA/zaD26uLda
IFzlTNsjo2558GmNUhM9FRMRnfwpe0AQ2rO09BjZfEv/WfKv2LsjlRDYNA821TCMRcTX5fUqEYPR
iyJInPlb/7sIklK+Tvpe9l9x7/cxP1DEeN5J+DH14qVosvKpHiw+U1nPa03oHw8GpDwUhws4zKy4
OD5KlJz4Oc/f/8c/oj9ne9vhZv6zXYu749dmMidwUZplUiPaaahStcPYgo/bzfUdXubbZlq8izM7
ma+fwQuMDxcmrLtfDecAawmk6m/JKSjMk46MlI6NZoyVDbScVnNo+NY8TNdVtJmFZEqd0W4O76Ed
jAD88G6zkD0HitCKCsAEp6qeZWeWlymdJcxEEYUIyS+XaPOmFtqAD+Sv2xCVI6m9vTdGPfBe4fan
lRo2PRLkzfQw438u6UsH3J2QscgT+Mh6RPxUTcQyUZjAotgGetdTPWhD7plInVK3Chm2VpAyClwR
xLL9bZrztaHrQfriEMrUjR4T4wdC/AO5G0VPAYqzyRfmZ7Xq3leDOtZHeXBHJM/jHEc7y6LvSkKB
rt2JWnnbMTaQqmybXd0=
`protect end_protected
