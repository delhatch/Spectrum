��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�XI�oq����P�^�
�{�7��/P�`n�1���Em4>߈D���_`VQ≃�E��=� 3Y��]��$��@���ޣM��s�X�U4���>6��D"n�G��A�H��YC39�N�ܻ�}�F�D� [�"��Sl�c�䪧Q�~���}��v�Ù�{~�z�	�vt�``#��\�nv}���+=�	o��Z��ʃ����_��xQp���M%����V%=��g�ϻ��q���̽ՋS�T��c���8HL ͫ�hķ6��'�h	a�2~h:cE�w��	1QmSy���KF���	�`-�Ȥ!��7�Rԏ3	t*���һ�)5��6#.�C��WkK-��eyxsEb�ӯ�O���f�5jهTڛ�a�Z�L�K�C������vD���-41�Y�1^���Y�U'q�<��Дΐ��'��y֕�� ��ӧ�:����Ո�W������ҽ�Y���Re���Ԃ��O���z��U؝���r.������b�&�Dzg[#�|��U���h��
1�8���7'[��|~I�����)#��7�J�<<�ÍgF��P��]%�d��ZK"��@?8�̓<N/D��v���9a�%)$ZTZ)4Kީ�9*兇y���!�p�̞>}�I�́F�4<~��O-/Xg�X>$��D"��1���~X44$�.��P;�x�5{�O|[���:��C�z�
�dc�G���I�K���?��@?��K\��0*��LkZ�5���`Wc�(n��]�@���DQ�N1�X�ƙ�m?HH���xz�aWQc��o��b�^f5yϽa��5@��&J��ǎ^��?u?�WEF�� ��nk�.z��V�:����i���[V<��u�_�l��?ŀ317�S�p����J������¸T�ͫ_aR� ��?�Y�����{�(�A������,|k>�a*(���{mrҿS�,��$A�K�B0��8B\�O�i0h�䣋��{h`��O2,�g�4*@+"�B?�8�G6lv�����$"yy{�J���
�db�,�,��洬6�����\�
�ʨ>��9G~�
�)�������-��xA��\|�\���5&��~���	zg��|�a��Tь���Х0/���C6/��0�c5�����>�����9v�����qI�1}!�t��[��&5њ�#ø`��ո��n�������D�l�N�ΞoF�2�Z�$1��S�&+��~ف��~G�'�d`�m�f[��*�r�'�^��g��Ե���+�m��z�(y�����=���j�17:7DB6�~xB�@�&�[""q��J�@!�H��˖���%��E޲�@V�(�)�!� m*�YU�}	���U�~����!��/~����">��
|���#=�L^R�++���Jw��)��\������t�N��ܖ��!d�E'����CI	д�+v��I�u�> ���'k�����tۋ��c�i�q'�ZD	��ү9��3=��'L�|���W� 骷4f$���<"�m	Dj0�r������[�5��Q���b�xaS������ղI�75A?�h��7�;��iI��
�̅U�`R��Yպ�|�Sa��]	rx����A$p���!5�L#��?�#g����R5���D�ۆ�X_�;IM~�Va�r�^Y<xpa��V��e���)$��T��G�A�o[���Z ۠�ά��̤]%&�)��]
K��m��o�}l�Ԣ�oK�۪�`��|�ʅ���!��-�Kf9��D1-s�}����=}K�b��5z��g���cJ�]lp�����|�m!�$\��@��roa/pxB�lk�"D�+M���)�����M�"�2U5����K���ez��tk1�K�^����K�q��բ�,7Կ8����Y�SGP���&��\AZw�}�ÂewQ��K�ޤR�K�`ݳ)����
G���(S���
#a�ģ[�:�{H)].u�ڇȒV�k���ǿ����o�7��� �T,����!]�7V�D�y9N��zӯ���h�J`���N;��|� ��������1<~�Ӣ1���Z
�������){L�A���Z'y$�<3z��;���3j��7����!�р��mѷc��'�{/�9����VJn�k@�O��_����E�Aѓ�x(MK�_��b^k(6rcY�Q*�6B�=��wqW�`|�Dx�co f�� �E�uMC{Lg��~��Nm��jP|K�쎁Ο�0�*3�K��=fL��[�l�Ƅ0���\��ҽ�=\�[�-;p�>��-B���@VH��ڴs�dw���K��}q�V�jE�M`����g��-�TC���T$��4��r���b�b�<U�.�.���L밲��'*N ?8x�A��/X����q&����Z�mM*)�Ō�:��N}�hw�����11$^�Tϭ�t��^��5�:�.Kْr1c�P1!���R�X����O^�G���c�d�x�d6ͺ�ɗ;p�t���qǃ����US.dڜ,F~���7\g�����t�lSL�s'���i��<A���9,�W �@�=�3���'+��f���#E�U��:�c"������+-:^����)m�,P$�}\Ѥ����߻��ޙ��hE,�Ʃav$�� PO1�l��.iC �]�dKu��׏ʾ�U�@W��s�2=� w���=UQ�1Jb��<\���¶2�!R�3�J!Tg_-����I)m�a'�1F��\/��x�Z�yv���o]����E�A���r�����&ϝ\aT��Pp��L�9N��R*o��u�U.�ѹ�?]Qɥ�1�O̎�eR5ķ���l��4��}���ԯd���#^Ҵ���ⰢO�/�2Kw���"FN=	������K���_r��4:���dY�-7S��"X��R�t�iC�c��w��y�_�w�{D��15�����=*��}ݯy���_�%�l@��1�[��ǡ��'��
��&s�>[ݏ	n�o`������� �8��MR�k�B����X�?2R��B�z�|��:���#���B2���aR֯"����}�|��8{����6�
d�������;���ĎX�5slݚI�j�����<ZVҸݟ-̎�b :,���������"֩ �.�<���B~*4}�DAex�Jq��	W"�߭�E��
ώP�t��"y
4�`ê1B����S��ʤ>��聴�~��%�b�%ɭ^��B-_	����
�Yc�Hɖ�2yN궹�U��(,
�sR�Xc�ǻ��м�M׵9l쎮��VHؚh퓇g��e���;!$���;��Yp
��Y�]��W��u�䣸���˚v>+�������$�l5���'�Q��9�����HSӃ�x�!)���{I���췩��O+��RX���${.����P�=�����t�W-��%@���oZ���fT�O�}	o�s4f�T|���	��`:l"au���	�w����O���f�ls����͡a&��{M�t��>�t�}�"S��G����Y�z�d��w'�6���UHC���c�[�s��V��w~҂����j��!�2��a�bq���u��}��E�W}���}�h�J_��"j�� Kw��t����Θ��Ulq�u����:A������i/Z^�j�fh�y���;�M��7�q�ds��M��h��Q_��W7y@�Ǆ{Q���t�_o�%hif)G:z5���Q��/oqkp�ZTa��1��q��U��� �K�S��5e7�ש�R�w�;A%�^�;8�3m�2" n�ѩh�Qj�`^���k�Iʛ�Tz&d���
(;�&cM�x[�f���O��8}���~z�U�#e�7g�W�8�y����RZ��ZQw��1gw�H��+/TW�ž��Kt0?cr�T}E�����'��f������_�o��1�7�s�"��)�A�<��hf���%T��d�p|2����)�����C��#�#�K���
�H+6���⍵3�:+�-�פ�'�}5�s���Z9`�g5��D�Bj^��‑|�����s8�Z�pVN&�='��EZ������@��ͳ��2�ed#���h�\�֓F�ϫB\�Y$�,e�%_><?!Vc#	dlo�nj���x3"".���e�#�$�uhh�0R���O.r8��&����`[���J�Zi��k���$m��2ˎMG��Ajϭ;�n�V7��OeJ��RQ��|MY`ޫ5���/��&^ �����V��w#�"�8���9�=��o<���`<�j<꽈tc֦�����Bˉ��@�̖ Y��@c����]����lX}����\b��<�/J�'@�z�
T���ٍ�u�c}��8����I����>`w��v�fZ�m�;���Wf�f��_�������si�y���J����V�s�
���ߠG'��K��"y�:ң�7q����[hR>�.���	r�����g�y�HL��C<r��UͩUO&`�fq�x�������%;_��Ӫp�F|�p�%�����Ɣ�X]�����װ%m�-;G  ���\����:�T ������ :|�^�3�Z�����	���?��$]8r{5ٮs�L�ۣ�dx6��H8D@��ضԽ'p�v�Y���a��q�"�@>pv�ڪ��6���8�}tBd-� ��R=v�] �S�W��'�,`FA�a�"�|�N.�@g�Ai�� ���<���K>y��wZw�x��:խ�N���R�~�9(b;�/��+$�1��2��<2�.rR����ծ+�&]Y�0h���Z�<�9�+��U-my� �a��C�����$M�+r����h�H1*��Z !TJ�2$��Ա'*e��-bO���U��9�Qx�6���<�7�o��X����xC'�`����Wߗ�p0����ԏ��U�AwG��)��f���'�k�"6ß[��̛:_V��j�ķ��l��+���)����`����L'�;�퐶�i�2��������$�P�3�E?�B|�~� �O}qP�OH�g6�s�rՏ�:o�:����7T�%.o��h�ј�g��Y�WF�r2RM{�a�>B�e��B��w������/�`r���l�9&�M��R@w�3�1@[|0�D4�]NS��Xq\�	�#Fe=_7�<x��33��<;&�YL���yf$�yj�qZ��ɾ�8B��@�#��=:N�5�_����!������<�WT�:,>y.��(~�V�~ ��+yy��YÒ�6rqT�+K���`��!�iO�7���&X}|PZh��>����(���o~�O=���W6�}^`�7"�_>�6Q_��i?� K�g���9��I��`�������&��n���~�w��\�0>~��Ff�?��8l���S��e��f�(�T��F؏���>0S��4��P+��_��Yl!�1Ji��q09C��K����x���'�u����)#�d���Mwt,��i9L��m#
�u�Y���<���ԫ�L81퀿���B��J��MmW p�T������	?NΒ>G��l���Rf3s�yv�@"�wy�����}���u�)�-�@���=G�+���h�c���t�n�����˙��9�E�x��.y�g�T"��WL����V	r�Z&!��X�; �!���1�[�8z��q�s�#��eM�lЃ�U���5
P-syt /�۴z����[�\7'�癸�e�}��Bs#�|�`�Q�K�r�,A��Pm8�{��ރv֫�]���=Y>K�@:-��8�/Ps��.��Ɍ�g�"�w�� zԍ��O�**�ESǚ5
�ݯ���e)�n>����W��O"܌�U�EG��U�G��wf���"�1�@N���C����QG��0���Z�>Y��fOL��H��j�5���0K�g�@Z�O�9q1����b{�4�ۈwH@.�o¥7�6s�J��s>N�%o^���!��sT��|a����K��|�\�X�]�:VЃ\u�B��f#z���/�{���Ŧ�b͇<St����d�]~�QҚ�{�,��=O��@�D�ۼ	2-�b�[Q'wv4���ђ*�<����γ��RL�;I�޻���c��[NL�FRY��\G�;H�gҩ:�� ��)�4�d��얈���x~�?�����Kg���F��C a����/H��'EGpWO/'r����}�3<Ox5��CV02�!s0��hs�� N>� f�%���|��µbh�g��j�ϻڲ����L�#w}o�nG�޸\��@����D]�ɠ���BO��4E�82�I.��M��!m�z��ǭj�h�oժG����-aʞ۾4�����b���E�%�?D��;��ÂٮBa6;Sr2A�����!c��{�@�0��<�*�U���H�)�P�|N�O��
;]T��p�s0���9��ӑpY��Vd���)�)�T�0������ߢx�`�s�1z�.3n�R6��R��C�hQ�9�R5�|���ݗ�R-��IU�[�.{7Y��z�bE�{��߫+�	[u��U�����e>���*��
q����$���ͫ>��خ^���#1��咄`5l��]tʒ��B5���D�U`��ū�P�^@S�Ah�9��v@ �X�~(R�p1�X�)G�p:b<������C
Ħ_>ki"{��9�n��jb��c[��|�����i|\S|&��C:�K��:��s���ulF�Aq��S=����E�3����!h�L��YOOgDZi�_jp���U�!Y�����7�萉~-�d�J����������
)�dv�8�ϥtQ��j�߭Y�6_h�����"5{�g$3-kʦ�����nS=��������c�KY�Tz�- N!���C�ӱxA�ey-�<%�x"N6�E����#3LDY-��s�G��r缿O9���c ��(]�6d���k޾^)�@�o`be_ţȿ�w�<��~�!���~�}�^�rЫ���KR��U_���?E����'"�k.!��R��2�f8���:�7���� |g�nrA@�ݫS��� ����޹I�_�aO����6!$~�i{5�$5��T���L�ںLL�_�ug�ƙ">����hՕ�z��?��V��;�����o�dnu�B��)h�)���C���\��'>ߪ�@N`v�"B�0�p' ��P\�-�] ���>r��9d�"|IV3<�_�5q�L�n�#�V�,F�{-1Ћ��X�����u<��4_��0!���,&535$�22ӏ B��忞��[��Êy�e*u���M�"�ǲD�����ud�oa��	^%��i[��De�X�*y
F40f��8z,Nn�/�t�繟�i�/]c�	�B � ���=��^�q1�������n���Xl�%^R��$��q����E_A���NlU���M>�^��IAߕU�<>n��_��DP���+�r���B9I!��ڡC��X4$�a�GK7�~�ު�2`�:e��@��5�ķ�S�����!/Єj �ݴ�c�(�"k��!e�-S��9�c����X�hS{���W��D�]��U�p�D�H)�(�1����?fdX�ẁ݄��f�&�И�sT]���m��� �i��BZ�z��;��> ����`��t�ȇ�f����P���6��9A�"�a��O�/�sr��⡍<�\���3��ɬ��9�?�롰�HW2S�Ǎ�0y'�,m����>8���y�e��
f�<�&Z**���t�z����C$�u��̽���+T�Wr2��� �S�͊>Y���极�ᮒ�Uߒ�o�M�NmDb��'(�$9�=��
J�U�˳[���������K/g�h�"�P���Y��S7z���+@�6i����J�����A���%V�~7Rh�`���gj��@��k^$�R�+�����1zӃ ��**�$��c��v���_��@�h�c�wF"y���>�t��Be-:����E��N���hP�)C��;�P�\�S5G��y��2s�P���Ղ��wg��'�"]҆qS�iW��C��W��mp�?T�]}|j�����&�/�����Q I�N/g��+�4C����yH���;��8� ���k׏kT#D�1L?'��U�7���J�% ���H���f���k-���1�i8<h{�޼�c_��\�N��d�д���z2��N��$cE��9��.s�	�AH�����3lNp�?��J�$�ޙvN螊�ؒ!B�Ɯ�e�s��`�D�B��I@�Bx��_��"���	���ѷ{��t��<*i5�?:�J��+��q����Ѽ��4�38�+.N�J�Ymg�����p��Hxn��ͺ;�����T�[ų�f�Z��|�߀����b{���g��z�;��u�ᝰ�g��Ւʱ��Y|�.���Ծ[N2��&��0�b�}3�l�= �1̞�!�WJ��޴�¯�ßQ�Qk�YDG7C�,�K+������`i�}<���)W�aX��5q-��w�r���P��`��r���[��oxf��i(�j#������ ";���a(eԜe!B7ޣ1�\6�q�Y��&�|��[�uj<;�2r9�_�����b��qs5��&g\�j���s" ����JjW��u�945W�̫u.0s��	j	RB�`��Tc��$=5��SC�`4�%f7`�=��G�á���U������c�gF��00X(���.��h��a'�����H����������=�S(2	c%�{�N�E$�$�K9㗋R�hʀ��4�V�֜�pd�#U�K��+������9���<ԄL�$�JQ�ʙ6z�U{�񪧡�kt�SJ�f��A��쳡{R:d������U�/�>t�v-3� M�̕�tBx͗��/��1�6���+	gq`�4�{��Z;Yw}ښ>�(��$�U�M��8E�9�⢛�r\8�?f��M6)�}����̔ R�^�Xs\�kDþ\����'B	�^��F/�Ϟ�_rp�(SO)�����^�֓��c{�kg�I�]50_�3��@&D�A!��lpk����a���2�~ڜê�W
���'��o�L���-`��T8�dB�q�RQҚ�zـ� wH1g�7Lv)a�:� x��G�S%��
8�/<īA[������֎\�������w7-�lSh�l�����8�2�o���F�m��3<���3� ׌�tm�կ����Uw�|f�m�Vk3˪u x(�����,���B1�a ݻ�w�9�%�!��y�`,w�aqJ�]�^|�#G�ŧ,@��c��k��~�Ԥ8d4��&�tx��`��<z�#|"89�� �n�G�gj�b�_��R��(���%L�1OT3�rPjG�҃�{���to ]H&GͭP[X�y+R�됟�=s'��!D�\ȠM�[�Wˣc��Y��r����ũ)��+��@%8��f=�:�T�N-�Z��?H��	��6�m���X�^�k�6eC�/=|^(\��T8΋�&�JAj������N�?"ˡs��0=�'����oRV������TX��\��������T�[Y��cb��4��P��Ԥ9�ي�Rƴ�e��+�8�h32%�Wء�G��q�9��M�����;�1¤���}�������s�eWզB�z�����I��s��$v0��7qnj!�	�ᰯ[`#p���'J�eo"Y&���}�pި=3�K:,(�Kd큖e\�']�� �,���Nc�w5�C�׵��{*&�{���:�\�̰	��\K0���p}��b��q}lTI������^�%�V
�����A�L-ժ|�]��0�F=pm�y4A�`ל�N��}|I�p�(�LG�慱��~�u�U���'&�H�5�L&gʍ�D@%��S.�&������>�!"�����v Y����6<-���r�̍>����#_x���	`�ԓ+[('\�����	*�I��𚘟���2;jaWdg�^n��{eSꜴ S=��	��)�_1�eeӁx�3��Nm��dvZGM����K��	�|�O?c�vG풮Fu�Ndf-���)��?�|�	�f�:g:I�9e����PY� 0[��R���*s.r06�8�;�6�]v��NLG���v��G9TS��D����{���)��|y�L�����$�97öG� >����O�8���f��ip�>R�X�-�r���|��#q>�a�)�R+)R�ˬ�B�QxP�+�aĶ\Q�l�JSuT�ɐF���e