��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X��q�{.]V���W>�R'=$��xr0]�i"(�����<{\�����������w�:�q�8W�I��o��,�9�g*�R�O����J��A8=_��UHbx�1r���[�YV%Z�)��Q�4ΏYȊ�#i�*�D)��s�:ˇ����"�&���-���'#��^��(��U|p[�=L�������E�b0e�p�1�ɦ�>��I��۱0���z"�ɂ��S����2�B�f���a2ic[�\�2;%(;�ꈂ!�K�)@����+n��c�~�Q\���B,g�d����i�a�(�<�6(�	3���w(�Z4�p^�m��neIB�{\�ü��`㟪	��!m������xИ�l)����=��c\�)�j��|'��	*��!�'�����k�8�c4���N6!*� ���k�����}b��xpuľNuJ���;��� ��D�ɋ���Xλ~NT]8��˽wI���ݼ�����Co�� ?*�ȍB3S��r`)sŲ�)wid���~�[�P��9��%���3AFw3�<�𹻇k�W��`�zk�s��NM$_��g�k�9�8iX\�,��f�Nd��o�۷4y[��1�Q���9���	&Q�!A���*�/��]uK����ܹz�q̄�����)-#��0�� ����uEG
��9S+QΥi��q;ңK���"o1z>����Z� ������
��=�@�Wi�y<���W�iv�E�ʽ���;�G��4�J^KY��'�i9_N��H�O����כ�3�n��E�"����u=��n�4���xu�
@��ˡPsX_S7٬I�7y�Ye<ºS#XJ�������>]�k�r\V����lx��j�4���"Ni�A��vzl r�䇔����t;�ǙV����d4h�H�2X�u�����wa�7t�WY�_�]fL��t���U<�{��e�
��4jv'sL�����R�'���%�ɝZ�~��5>���!j�����9ɺ�&,���x�
��tdR�u�m8�������ρ���a�f����8��}J4� ���T��s�.nV��Nt��d7E�$��i��!�+��ѷnW�## (@�W����Պ!�Ԡ)H�7m��t��CFA7�ñ��o�zE���0�Ү��Cp)Op����O�oW�3��KA�㫼	5��G��>�"�� �0��A�-���4�r*[��,p��=i�@�.9�����ڇꐎZk��-�A��֪?���7��� �v�����-��6=��r2׍#��Íx&K�ݎY�U�����B�'}���WUs3�M轁�fN�ڑf�$W�tZ{=�iȘ����
�է)3#�<#����nK�^��zs�N���W��Lﾧʧd���O0�Q�Ա����I�����s����I��W�d��,~t����$��ȞO�L�F��<�ƀ�j��p�;��h�輭L���1$��Hџs���(R�k��+Z!d]�%�x�~mw���KT��w��E�g�,���r��;�`:F�U�Y)�CFo䂵'��'����F�P������aS��WO�pm��s0�\�+�a�߉5�,��T�:�}~�G"�:1���AUЖ�v��vs]�`�J�6�H��؊_WF�J�<AI��t�u?H|��^��X]P���N[���\ɽl�� �QegWS��m��4m�kAN����'�әW�j�������u�����C�2��0�\0��ٛ��X��7������}t�L�Q�%%��Ғ�6k����bO2�H�}�^ П���s��{����5��HRkO��I����,HHZŏ�_�S��AM��{Z&�4�{V���-�ŬpW��pE�iE�7R{�b��͘6�6��cO���7�1��ҩsy[����g$X$ջ`�j���*��Ǝc��@�-�2T��O��W'1b�B/�Ǜ+�c����E����	M��HB�#I=2c,��N͸��xDR-�.����,m�#�p���9��ś�0�P̔J���(�Fp�%:,�)oL�i�b�)����4�_�#1=Tu��[�+9�u[:"����qj�-���d���ٖ��Y�<�fM�w�k���ѳ[@��&':J���������0���w��Ћ���4��G��^'����3E��߮���^��*��M??��g�uO�M�]?�g7Hu:�;A�hYO�w^=����ʥv�/��緊!]|��U`���6�hQ�W�)}̯p�*�(����>$!cAk;��Xk����}~�����1���'�T5	���݃n1�@���w��A���9�E��`�������0H �)���Y��<[����4a�=!��&�r���>������
�1�Jv���
����������@�eW
��h����!Yr�MHR���5NkEW7A��rhd4U0���*�gG?D��=I��V�c?=D�Q[�&��-��H��J��CmkC���&�J�6��������ǺgrxF��Y�yXVuH�=�#U�
mp!,@��V���)��)BkTSJf	�G�Lw����<N<� ��� �o��,e�a8�p�ڔ����[l��y)��7N��_%�/o�3;���6�dP�j��Wnn�[� Չ�O��M*��G3^��%"a	���P�p�<�gҎǌv��\Gu:k�@4�����\yݔ.����j1���F�(�sއaU�2����bV��ި��<�Ä�u��y �Gg�Ps9�_�Yp-�J}#���_s��7w����3{!:�	�d�������m��I�BK#�[y���_6���
/���1��ȏ]�/�<E�_.!���B���
�6��`�q�@p����S��*�dM],'_P���lJ?6̏��s�������YܠFD��V�=d�hzP+	�{Vvr�|�II�� j=�R�F3,(X�3�|����K�����=o��,�1���T�t
@'����=͏�UXG6����G���8� {G�MN��>J���{�A@~�����f&�t$T�Ur��?2+�l�b"Ё��3�C	��ℭ�]�&p��L����kA��=F�4c~-,Q�)�yOV[���cC@�}_�.T�?z@<��-gd�>�1"#���D��������?D$F���	VN��mM�d��rr�Xu[y��pP�9 ib��LUJ�������'um�؝�纃�O�n駤���2PɆn3b�6�X_݌�
S��$��j�KBazyAItּ���~�ZP_͎�S쵒�U=A������*�^.zC_����?�r��a��]�t�+�,rg
6X�LtX��byJ����%�-j1L��N�}��[?`��׻&y
��6r���+dD�>n�V�SB臈�oD�jC�,�R��/kJu� aѻ����!�?h�d�=�v�.B����y8ghu
Έ="��a���p����F�@����rit��S;`�K�&@���l,���nqK|H�:~�Hze-��❗|e�,��;��#W��ݡ3?&k����7�R��I��-iE1�3F��Wg���~�г�s&N�;�+���V>L0Q���|�X�;دa��M"w���q��)[ZF��*���,Ĉ�t��S*B��?P��![�mc^q� K���` �ڄ����ǻ&LQp������Nn��H�	���~q�Z=��E��V�zŧ4�E�ZD�mQ�	.mB�U���'!��\&
7�q�=&��P���l�F��9H&N s{VڒX�����ƣ,̷�ee��J/�3aP�=�#(<��7����d�fR9�n~J��[+�&�ܯu�Kug�yIh��&�f��!��n��x_�T*��㓢L��>F
ɑ=���C�K�3�1��đ�&�A��	���Ȩ�� <@ dՂ�b�>9��8�嘮8��;I��n��!�UQ�T�U,~!��SS��=܉�>!�m�
E?ׅK��������J}�l�	�#��Z�7�+z�}xƯ�/?���/W?���
4��2ʞ��
~����G~�Aφ1��usj�����u�G��h�W>��Xhy�[y�^�����5���.8[���Jo���߀Ny9���t:\e4��B5.�<���׏q�����7p,pS���<{[3=��2��>���9J�d4L�{�^�r	T�|���ē�Q�y�s�h�8�å��ʿ;81�r��%�S�h�C����J?^�$�ݰ7��`iUJ�6\~�
��`:���2��V��� ����0Ҥ1�G��w�O�byf�op�o� J��P>3V�=�����}v�D�KҴXZ�����%�_����O����)�Wg�]%��ҙ࠳��mb�%��J>��6�`\��ѹ$���+Lf����<�Ñ�7�=%��`o/�Mw�7U��t]A���w�E��6���[�w�##M���z�׼o��Ճ0剓�6k��Q�y+8�%Ӗ���ړ�Z��Ö��$�4K����S��IJ9�\��:Y�1��b��;'j�,�Ѓ�������@3�}Y��y�៾��cףK�Ϻ�D���v���"�N	/�|M�Թ�4��D@�^�/	޾�S'��Z�J���\*��;5��B�����M��_V��kOv�}+@�;<��걊�8ɨ6���^<�R8����#�yn�!�,��E.�����0��H��k�����4��tV5!���~�@���{�d��Ӿ)Xn����X4\�G����d����PR��c]h�3�X&�����n�fT��X�	�h����ï���>�<�+y�s�oB�;V��ڝ�59p/����� �5�(`e���[�2 ��%S!����� ���q��<�o;�y���Rk�C�C����[E��X�����k(+���t��Q��2qfKy�u�t6��e��g����|iܝ��V�F�#9�Acb�D_,�*:	���G$ٱ�BE5|Яe.��{�X���^э��"���~�n��(L���no?�-�uU=Y����u���Y:�p�=���=o��F���7N���q��=��WX&ׁ�3�5���9�YC5�_�!�����9L�?Y�>nG�(����_��SJ��~� �L�V�G� �W�B��J���-�7`�.�3�/��*�H�J�u�=�:	c�O��*�Ae�����Iu&k���u�"��--�8`���L#�I!�U�\K#$<�B�YSʴ�2XX���e