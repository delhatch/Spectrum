��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X�@z�|�Z
���XL/Q,�"`�;G9���;���7��y��r{v���\y�.::ht�lE���R0��i5����16V��(%� fx�N֖��c�8jK�SuP� R1�:%�тT�7�?;�U��@f?Tdr����X���8��:xc�J�ilG�Ҝ�US.�EP�U&�Ra�[�	p��
�5��n���=h7�J�J%h���n=9���&�t��"����r@��'ߊ� ��K#s۰����f�	|K��!����N��"J��9��i���^���VuԣW��uXp�&Fh%&��C"_5�N\�E��i�T�<D(��5�*�+|0*�L���������w���K�k�ܕ�`v?~0��4�"��X�\كB�6�~HI��E�/�G���a�z��n(J�?�x3�ML_���m���r��ڲ���B��c�'��B���%!b =S2	���<��}��.��#�`��0�թk3n�����Z��P�Q�+t�=L��<[I��aw���p뿗��;U�D�ܑ.y2i�j�`,�}1����%TFn�eyuO�}�K�Z��3 j��ŀ�!�Ӫ����$�E~��[�ʈ����ͮ@���{xץ� h��1=���9��f�|��2GC�[D8�Ǧ������hb^���S�xZp�6�'�\�$���R>��`7�����X�`&E��k"T�ّ,3x4B�(Q�13+�-����ć�Qʓ��w�ӌǚ�U!�8 �ǔ6e+���'ۗ��#r�)(~:������ݑ�G-5��t���p�����9Q����T�x{B���vͷ�c�U��OkeG^����<v�If��n���m���ck
N(k�#��D�<ި�$']fl����|~�� 
Vd��\d,�����mÌ���:�Q�������|/�d��|�P�f9r�/vϐ��+�`<K#�S>�Q�hc�sD�^@_�>�d]-���B& $�Oq�	 �_Pu��k��9a�6��9�䅺(K��G�v�z�{I�Kg}�v�s�?�(ae��]��D��P����Gi:��^ �����S=��?q{r���C�!�BA;k��b��:�i*�T�Њ�����:ǯ������@�"р���D�
5M�kEj��[6=ͥXѢ.a�Qx��͢p��Y{�mC�\�P}]���gӜ5
&����v5xh�qR"t$��%F��؍_.DC1)�3�����#48����K9����f�sMYF(�>&_�/��|���%�-cV4�ŕGŊ)[��@ˑ�{?�),�x�uz
J��а�p5| ����|����kNmḻSO*�9kej�l�nc^�; t$鄺�ս�������H��g:�_ ��-5�l�)�>�͏�&�����v��C8�t���F�t<8��d�
����).0�&D{���Zm]d�2�mCg>>��Ң�#l�CvΑ���v�Ȉ��j���,�*�B���}�t�j�)<&[��^J8T������e��gsL�Q��:�7�x�X��]wA�c��~��gw��X�D�z�l�qN5fl���~��e�gk�����Z�Yo���⬴�iὬ��J9b���@ӛ�*I���J����l��HΚ{	7�=�� -���-�'����	�17���oǀ���r���6���IN��n��1��/�4(�Ȥk��T������a�� S�u,���1�7�������(���[���`��*���8�:Dθ�ki�ŷ�	���Df����$XXE�,�}s�#�g�+s�9�%j#^���Jo��k���#Fo����GRw�����[�1'E���i =�FUۘ��܎}@`�j\��,��uu�g�>�������F�t�h5�������p�*�}c�����c�?�x-����Sz�[�A�RQ�z	��@+S������g�ÊUAE����|��}Z���x�q��v��M=���~\P����i(�X�~IQ*��ɿ��°7
d���!Nl��vn/���K-i����a����M!.ZZ��p��a��j�Z�t�ה�Dr��I:�m�/d��g��k��yu�3W�\kq՞�t�m��7�U������'v�D���,1QJqGz!��\h�Oue���Z֛Ǻ}��Ż�}TǧM;��y7$�A��� G�>N�2�����Z�k<fS��J�~�l�g�y��?�Wb:�X�[�B�M^r؍w�U8�'�> v��@��/e�e����� ��{FQg-m���uA�ʶ��9A��!�q�1��N�T�02T���2��G�D1Xj��;="�O�h��QE��5���M�M�q{Ck�c� ��S�F�o��Z�Byt_�n|{CQY�*Mud�h� ����\'��fTm �xiq/67�r}37�^�7sR"x���\�2�K�;v�-��L�r�����d��Ây����a2;�듕�:շ����a��Pf�-[����k)�g,��x�@�S�?��9����F�h��1dI��U�&��~��;�ڏ*+���L��t�����\�������_�;��9�UZ8���Y�j�g�I�iH:�;�d�`|���r����*Æ\3�g��A9u{j�@����v�4ֿ��M܄����e�{�� W�w�m�$�^ؘ�vȣL����o"DUX�
%.n[��[�VCx���,_�As�&5a�c~�]J]��[��ݹ��UQ�L�:�`�(�l!�^$Y��=�U�NE�j/�yU�  d��lޕar��1`��Kk}�n6/Pv�k2���P �ϳ%4����a�l1�nr�#�H�T >fCE�kQ��S6f=0������5\���4��ճ�D��)��m'�9�N�x2(O������Ϫ�4� �E���z��˅L�=8�$;ꞽ~�(��!�cF3�>�_8��S��`a �p��=R���
�V/���fp�AľuZ^�؊@����e�ޠ!��d�YEX`���N
�&|�.��{XK�0�"�C²���3yIy ��y�������0
"�Y8�3��F1�H��L������B��[-y��Q�`�o0B[�|]�J�hc�+}�Qp�y��U�u����>f�ۉX)��>���Z���^c��B�����B�!���6K�^�H��� �(����%E��^߿�0�?�+�~��^������0U�R�J\�Ձ�a���k�Q��t��`5;����7��:�gP�Zy3C��J&F|`+Ȱ���kQ��;M\�C��C��Hw2�Qy No=�KL���+��P�ga�������o��M}[��tl=0&�؍X*�ɸ#�Q�X�(�8JgիR��5�O��
&�شFE���@�4=�[�WV��d!���̥Y�^��0�4��O�U�
n�}�9�`���]d]��k(���o�,��|")����I������Y���b�܀K;򂻎޹·K;5yp����p$�cױ ܝ��Yа�c�%C���FN���'L]!����&���_��j_!��g�I��q���i�[�y��'9;���B��Xő�5D���HV�𱋣�s�)