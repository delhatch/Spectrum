��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�Xuѳ����\�1�
֢��%)R���Zsbdɡg�C�E>�~�!��Q�g�a',�}@�jbWL??�dվqo�����
�>J�Q$2��v$���'�GK�GFKiSX6j���yB�c��e�p
��~-"�S�|jVޘք�T��R����Ly"}���j���P�j�S~C�|ER�*�=��s�H�#���bJ�������E�m8���t�&3��:��$�֕I ����W���#�mN�(8��c^I�k.d�v4��W�ڀ�]���TD{��ӕ��},��X>��)/��[�^�D7��}�*=37�i�3��6�f�!��-S����/�:�B�P%~X��
�1�7[Y/"����h'�Ѻ%0�2�M���i�G�)�,j^��r���)e��E�{�[2R�u��ٟ�-��*�;��p�����X)�%q����Q�.��5o���H���������f��Bds2�j�d�Q���+(*�P��]�Q<�@
�/�S����	B	�d�xH��I?3��N%v\f�� خa���Ǆ+�ѿ�y�}�#j�疫�Bb��<�>>�D�]KLS��}<N����!N<�VI�NPH}7�����U�|eL+���x����`��@aڨ��Vr��݈k�r�8���0��V��b��$H�DźyL>��飿��<��]�󢱝��NC'W�/�V�S���Pk�!�Fx�qD�v�ar�$Z����&�#6-�����DE�NQ�d9L51�g�Fa���lHQ`n��z?�H��o��p������z[��\�o<�y�� �I�VSyG����D7���w�S���	��x{�9n]�G��`��A��μ����_ޫ���Z�GmP�ʯ	� ���Жe'���:����&�"=o��̭;-���ȶϿ-�GD&����X�;���V��H5��I7��Y�	>_A��*��G��c��`��~��H�r�(w�rX����M�a@Pt���喺��"�{QǨSr��&0�$	܇/��ib�J>�y�b�K�_}Č�릮�NLdcbw �'�P���y9�e��B�FZZʋu\�x�B��!�ֻM�l�6�o](o�k��&�78��a0��l��!�������4�S}���G�<��ۡU���O�A�X<�qv,��2�x�����K��Vh+X�$;y�Rc���=����o ���FȰ���F��tqH��h�H3�n���
cusB�-��Z����@"��[�ls)�+�2p�+#O��~YI�'V
N��-��ۛe���{��eV�hs�B<(�7�����%��Q�a|�!Wzr���b���0Owt��x0q�HI�˒��:�t$A�� 7��5���rCCRN嚅1���G�|T\��>�z �@��Q���e�����6�!��F��X�s��>V�����0�%�7yXP�-	�=z�y��u�0ݿ���E��Q�_Z��ؽN����0����)zL�1�T8���m���K�y��J�V�c�_@h6��'�{�p:+���`���}�7��؏06�2���=�%���#̧�t�9�~YɌM��ނ�z`�7�k|XhȺ��j��v��%��K)n�OL#fG�@�rT�^w�>V�֤�"4Џ��xO��[����>/����7���w~h���,����q�fi�C�������1��_Hj La�;ok�,;�r�i�32 ��Z��?��2wQ:�)k*��?�����[L��W�g��1�ő���'�~C�J�d�/�i�t*�Nt�^�M���M�a�)�V�P��t�͝/K�p_�Mi|��4mO-�x`����G��Y�<|2��AȽش6үz�%dGwHC���m#Vr�d0��'�4x�O���,��?_����J��;ׁ7�"�����nr�����I�k��t�z�[���V�R��O-'��^S�}�������7�8�NW4�8:��7g�7o��~5�޺��j�*/઒7�����HQ�f�<���^ō�����F8�Ó;70 ��5E��0.�;�]F�p���G:.�5�ek�N�Ęat�1�)Pz�5XLP���٬�����R�r;	��a62{�Տ��3��L6�������(�	K^������c���y�1FM���ѓ�gE��[v�$�ئ0@eE��I���.�4D��0Jp_���T���Z�o9А�����ʦ{���å�g�Z0����f�Jk���F�O�M�	�=�����f��@���]��!�bK������c��݃��9�n8N9u_���U3�7X��4���-�w�Fm=&�	�;�����̬�q�+Jv&]L�
�o�z��O�䬬D���/A��f��#���~�>ݜ����v�LH-&1w�ȣ[�n��f�Tj��0�(�f�v�b��Q�V���M`�����9�����b�+�,�m�K����&�M6 �RПc�.6x�]�]kS��L��v��y��R=�y�D���a�p�n졓6�ٞ���M(8+��9q�t�-��S���$%vG6�@�O���Zj�;"��a� ��Dܽ.���&b��,�_<Hu������0������$��	���	�0�.|9����ޫ�u!q�
h�I��'?x��c���P�#3u_�ȕ�_%c�:6&�>���[��$�; &$���G/Z��7��&2��F�!:�^�X��2$,tv��F��z�H�0��2���f����O�db�ރ��d��<��Y�����.�m{�t�%��%��-⪫I3�K���=�J��zN��sfc�1����6��4@� ���*%�2��Eԡ��Y������J��O��3S�� ��iJ��:p$���N/�ӲD�]
2bgmQ0�4��}F|o�'L�`Z:G�f����ބ{��Y�Ԫh{�ST�)�9��s45�*j���:����G��ݵ���,d$x�#@Y�I�Z)��_����s{�^U�7s̲O�;�|��̣Pv�T���3�ԏ�	�X@�|nv�ϙ��K/b�����]iJ÷��۷�ϼ�����f����)��� au��JW��X2cT]o�N7��taJ'�)؊G$����_.�#��>ڽ.�k�����M�<Kgߝ����.�<ܰ�+�O�j�=�/����	�K=�3�þ��&Bw7�(O��rf��O�n�r精[��"�_z�c-� Fd��0~ ��H��s.M-�̚Q��#�*�l�愤ޜ�xv�oX���T<.*G�,sI�:z��W�ՉQ3ܷ~ۉ�G���ﶗ��%�!C7���&�.lVc�0\�j�c$�������{��wV�7hE0z,����j��!�l�BZt�H����jD���v��V]S���I �b|��8�,�]7��<��J'�}ft�dpvK����%������m,�|�[�	�v�qDrE���!�`qQ�EKc�b������~�{F�׃����>-1E�G`Mg�S�NX�D�X�8�oi����kD�B����]��ú�Gp�*d+H81�ن8t�Ps�5*6g�ʯ��������K�@*-�3��ep ht�Č�G~����I
�ʗr�HH���T��ݴFE"��'��e��w��92k/x;X�a��,�v���%ɄS1��=���~a"������U�5���&V�L,��ͅ�@��Yҷ�Q�+���{"�0��-Br">�E.�Ǥk�q& VU�;&�@e��ቘ�F��{De�XL�#�^�T��K#ZE�iJo��20�6nm�9���b��1���N�=*�w��������x$ u�H�<�<����J�)�ב~��l����[�&
u.�����$�����Xh5�|	��EmT���xZĈ�Qa��x�n����;�u
��cԟ���鹇ڞ5C��7�`���,�I �՝	��L~+����k��6nl7�j�=�a3�\.;n~��M��u�W��fqf����R����$HVxɹ����6�!y� d���,��4�#L�q�P���a�齶7o�q�u�s��ap���Ϝ�nb��;2$���)�g�Ȟa��O�������ES�![V��g��@�Ǵ��W�lD�E,Z�@��!������8�o�Q)�������sr�fJ̞jG�r�X���݆�<w0�+3�{9�l�cz�`]�oF|�A�����M�!`��4;�9����
�̓!�&/�}�Hq�^5�T��n�5m4l�}5�@�|:8�}|�S�7�/)[v�;��9��z����n�ad�V�R�]��4��O�+9�3�U���1���KD�	��}�l��-��i9#?;6z4��*�Hep�=h�Ls�C�6.�z,�x��B*:%.UP��7l��@��J���!	pD~�2�/t�M���������?�B���tI�D�M��gyDk�����<����379�.�ᣫ�*/�ؼ��'�C�h>6�@l�n�-2�����t$9u����7��)��x�b�Iv�g��lip;ϧIU�w-G?2^�0_����a�p�e�Gg���f������W 9t��E�py�;�v��eCKe=��c�_6D�:�Ӥ��4[W}/킱�<��Í�B�w~c��U�'&ހ���l-A��m�Jh�z���t,����n�n���Nw��TH�/1�4m�o����S` �i9|y5�[i����f���թ(�W�"B�?���ϼ Yo��y�i��F���5�q3�`��c��-����抙�g��So�B�@���19�Z)qz��
����\|h \���L��~�ؿX�]w �6 ���9Έ4�F�Owl(R���w6I4��a�F�L���*7Twp���_��!���~��`g��M���{��?!��'6	�q;�����V��{�$'��;�%1Շa���Pa���z+5T;S�Wa�Tr� �12�f)�ID�]a�� L�P	T�t������x�@�E����k���n���Y/�,!g�:�����{��:���#��w��0P͆oK���xc�ķf}�����e����M�)°�I$�C��GbS4\$�}}W�T`�S����$9e1W�/����/*����N`��j䯺�7"�b�E)��
��wY�4U86.��f&�J_*8�t�H�1�%��67��7 �3D�ц�~%���"��̜���G�BM3v�=(�d��@��,E\
'�a!,EB C���EY@�����E�I-���]j��#�Q7�L=�&���"�8��拍�H[�̈́�8���6��CF�7u�m����$Q��ꦉ
Y�GMp\�~��?U'����:-Oք��?H�m�hW��7Է����a*`�w&>Q̖���3�j�8XP����$�{�>��5��<�Xr���"��q�y3	q���q?x@
E��V�s!ʀب��୹L�dT�~8ޞMW��#��lr̩(*�Ks���A+y�|T��r�'�~�X��J{b��id�hF�0��sS.��=�;��бVapaG�#%I����(�sa����㻊��T ���Z!�
ٽ�{�&�/�$�6}2z,Zk[J�k�V�m�N��p��=���2>��DJ	�IF�>��97J��Ś$}}AJ��0��Ԭ0s -rA�@�����r��[���5�㏦"���ɷl��ܟ{m�W��&��3Ug�z�����VE~��k�a 'W��?18R� ��	�ހ�Ë+"�r���wȃ���.�va�0U�{��ۉF�
&̏��7�W�I����g�o�y~��x�o�m��cE��q����;֪�X&��|���HGͮ9.�e��q�V͑���0c��w!��y�����5i�r��`ȗR�1,���J|b�@�+J�6��O�����t�|������D^+/��j�r,8��7~m@ưf�E꜏�ըʗ=f���g�mof����g��S�OԨ\Ɨ~K��d	�w�wUe�&�[V^���r7��T��=ï����ҭm�2/���S��G5���V�F>�����y	��C4�b�O��(��#DҀ��.b 4�)���s7{��I/�T�����m��JD�����CT�UX�7����Ǭ%�R�>�2Ax��2B^|4@="������]���l%�8�ݑF�_�{KD���7&���4w�v�R�ӓ��&zb #���(8Dt@~�����Z�[��ϯ�v�잍�w�s�XzȠ�1�f����U�ԧ�m�z8�m���+/6i%�{�
5�̮��1r&�H��4��|�Zn�U���C�2SKG{hz�C��������Xw.^�Z��p�һO��@K�]7��:~�lv��*;ſ�B�k�iC`W�r�G�o?�F��@�V�mM3�UJ��+g���{��S�-GS��v̷c��L߁pv%��M������z��2c>7�ݰ7��x#��b�l��SWz��%D�͈�BZ
�_��wD�~c��E�dǃ2���֥Ll�Hk�3���{�8��O���"�
�M4��$��-��]�W�t��1��%�6���@e��2hL,5d��U0��f�e��K~Ɓ�N4:~h����
�l\��.�\�Y�\G���T^���1���*!KC4JZ	�arVu{QOn����t��TY%���u�ʎ��\�N��m � �ӓ�DI��|Z�Zkn�N��W%�j�eo����R�m�]nbH_��0�>'�Eֲ�@�b�x��%u����j�+P��y��u�(�}�[��d�+%�֞g��9�����N'�+h�Nk�Zq��8E��-%�D"�C׽�(qÔ�D�+��$�	�tO-��&?�q7���y�)��nK��Ԙ���F����?��P �x{��<3%�$�S��������xc�H8�>�a����l����OI��X.W*�04��_��eT+�rtj�7|/�*��̢��Gڴ���13y"/� $w���d_�J��٥�"X�b0&���%2=p�~δ	oMYH���I�y��V@��
+������@���Q���s?*HF뙬��mz��~D���w���,||��oj��� �!P�e��H�N�k25&�ා�P`n��/���3�TA�HTQ`�߃�~`�MxM���>��-a�ذʧ���&��u���d�(�l��#��m^����d*�;�
�r�.�B?�j��G�ב��j�ډ,g���.T`X�϶3��w��d��=��я�ɩê�J%k�Ҩ��H�U�����NYW��N_�n������.V(Q�q�+qd4y�H쳢v��q_������Ӟeo����[�*V4�jYFz�B`�1|�:t72�%Y��@%����} �=����a8X���/[���b���o�
R�|�Δ��xF0��;-��y��-���Ϭ��\[�Gڛ*��#�t���VZ������c�'�S���J}�Ҍ�q;W{�%��-�;K?�P�7��.���58OnJ��7]z?zu`�t��FF�jڮ��6^/~
���{��E�Գ��2�����I}��g��*�k��oMp��7Y��DN��KG��4�\���7��k����2��3 ��?�Hb4`�cΘ8������8e6*���]J�Akq�'6E��93k�?�"-���V��*��ڿ3����F�I�c��vj���W7��n��|�6��
Nc}=%�K�ZBS�Y_��pc8��q�Ƌ(	4� _�r�ͯθ���3-�����j�����\[$�B�K�1�Z�:.��R_�^H����W��6.r�K e�`M��J�G����o:��zq���Z�eP/�7b;:����_���_r��)�u�eG����Oe�s��ܬ�	3��[a�j�����8ɰ�ˀ��fp�~�~L�T�͓A�_�|(n�B�.t��~pHw0�V�_���������� �x���@���[��8\j?�	��� E}�JpȔ�'�&�b}(E:Z��J3�5�M�Y$�����׻<�r��W+�ݰ�W���9���Fn�"���[S�;�&��1Y����B�ӥ|[����H��j{��Oqô�7n�5-#�@
�����߲�H�á�V)��;ٕ��T���B�Y��պ�w����R��XJلQ�J�-��q'{���"ꪼ��E.�Z�&���
~�~�乾_{9���z-�w��A��)�\��Rr�,䯍|�D?��=��(Df��G�Mi-�fMz<r�V�{-�_Zn�-�G�s�c.��Er�'S\+�?�K���vl����6He