-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zIH1sKOhKWDSR0nIFWCYCAY4ZMJRTO6+as5cjz8tzONs8PQiKatgxqSfIXObzQzmYApfy8d/bYJH
+856zXiyUZiUkOMhaALpEP+v6Bc4V7QaoAWVEvcffWEVYbCufo3saaOFIyjsADnmUKGWaxk8tCKL
xAWinp8/fw+8KIW0Qfrkdav9qao8ItJnzircbM/y2Yr+NRgitB2uXfkWcYsjUfTs8FSK0kai/O6f
b8+jhKgfqUz5UNic4ejqHTie5YmV6R531VrY4eaCIXDuh+b5nMw39pmoNFStzezaqPagAN0yOAZF
uPU7RuZtFeMmEdJMuCBD+gIfucV8l2bvEwduqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
YwHv5/xY5di2mr6xHHGE3374ijGIp/x0UV/XN0R9rPU3u52GTPqCMBAMfuYwqCWLnNeiEJNNHTx4
qxRUzwT4hq5jZUMKRa7vpu5rxs+VhSl+KrzOYMRfnU4bmm9jFiPFD75pqQPimZ33p6c136JRReRF
pj4je04kuHuf4Tk4XUzsynZCJk2tNHawMI6Vtgiki2bJUxQDQ2G7tJciqeDS/R/cyKUKEXUutLCW
ts9X2RjZoat63ezDg2JVQtQZADvIRHCgPV40wnIo74VyV2NG1DKm/y2iSst/Du9vHPoLVZZ8Som0
Z4RnDCrv6gVN7Y2CINPIpmvwI40DL8QFX4z8lvutpLIeCUJ8vd4Bw9ndJML+bMzev0pprMN5MAbR
xx5EErwAvNz4TLOK9uqkA7n+kDF74zeIaQg9HZQGIOmWxWoc3kTAXDSA2Tf9wwcj5R6fQl4FS5dN
WuHiM+3qjse1BhDd7QhLcEhDnbMGcglWsBT4iYJRICmp7HwlB0nA+W3/ua1P6Sgzu+UgQPb4wiVt
P7h2VRVoz6Ut210gPfi6oV92Y4ZXi5bbZvr8vQONwM5mTx/X9RPrqTL3ENLgN28dK2Gn02e+Rx7j
AYtEdM76vxSvImTLkzAL8jwSoRd/9zt7EBcc8/bOpGxu9cFQWVZ5MCZ8jzNckdOn69xbc4ysftEj
GJu401/LxIIrmP00hS/A+u7RDjCaSuYAHPbcQbYuPHw9CwTArUb9eocZ78jmVInDfWH8qYzVlOFi
qIHMpqLvaCn7e0wpEd4Ywo/FKzLWVh1FWzAsPMM4CXgQVwd2lZ+d/1nYT2eTz8uueueKQnuCvivp
rPjGGOIj4MCLd5q/n9Gs30L9I/BEbxKsFeqN/I6sRZpiwVVEDoegQ6lkmkMDPAJJ7C7LAwUXyuZ8
hAkR+j2TR+hA17GZaMvU2afKIsF5t+aiGla3IchlS/250S42ux4Tygq9B28ho+A0Eis8QgOLoxQ1
gk11p4T6m6C2Ub5DthhksQeDsoqcarIJOsIW5y5Em5iZSwkxyj81dNek9miN0pudV8b7a/w48HvE
ifHnpQIu/qcdOdfUpUDzh8tQRp+m8vRekTpdtCUpuDYy6nu7TzRMp/HIbzgzLkMjuMlK+By6VbU1
CJsgDlH1Y18HTFWBbCgS0UxFd5xByDmDb6FRpMOjKFV1Lt521XgKguyO7N2nkWI7ePrmMw6SdRT1
jy1aw6+bdM/I3Iqm2C8ArRNefd8uGZggX9bbdAdVaa6htQPXLJef272p2u98V98rwMbTrBp23iHp
j5yjvSJbok06BDY/pn6VJNwEd4WB2ilVu+sMNnPwqf/cCloISAxVHyhTOLaNuhGXjBgv0sbfAdcq
rx7MTenWI9W9z47ZEWLztGXz6OmLSKlLuoVlFh7ddeCIQ5vXDGCPziuNvnQ5azfh4s6ZJCdle4kP
TjYqJ2BucohfCyoaKhROnsCsAF6yIroE30Ydq7Q7sYRNMTKhITOhpG0y86I90JLQdBlEtO9wskoO
3n8Dh3pMK7xP7+w436Y8BRwtw1tx6goQ/ZKfpgW2Dh4uOk9mH82YFqxl8bwz/3nVfMSiLNff4XWH
QjXlArahxc6BrjMuv5dTp7dyvOyrfWqMrFhaWb98EVcM7psJm0I4AgQOqbiakEJTpASv3Pb2cnNm
FPRls/3IgX+qWwpTCEii3w5sTrg3BwCy4BWHBSlv47MSjhtvoBjcZuR3tNvoADVZ4whs+F2yUeU+
GbwnG/m6iCY/lrC4I3AMEQy4FvtdNYR1NAxt9D4AHAsUvsSjpgXQHyAs3FqYxXPJPAnv2rRXrrS/
Q/49V3TTDUbQ+KgkZLBX6LcX8lJbvE/RTuAmsCzzMZuTli/W1HQMytBOsMjqpJzwnck9HMyWbbKH
ACRrFJJ43xWsLtTKAfsp5VwxUaSEvFeVLHkgZk+jttEOC9BQPpzZxXqZmBdBlcrGyZHwagsKbXEL
Twicim9bF1+va02uUA0eM+OiiQo71dyeHk/PqgCQDJ1EbD6wYYkZF9nXeqo665UUOUvZz5sEdnoe
uQtxwlbN0wU2bhvW8tuyNecKGOwOFqnjuKzM8lGIdodI+IdIvjbYqo83DMTekAxddNpr+BofyzGx
OtbYdmywjWlzihXM9GwIyHWMFBDGoxDXXx7lNd4k7e+9AMLQ4WcROEcIZ03FKtqOAeWsqTo104X2
XSYrBGNmSjklj8KDsmp8yGDelcXA0Zm8x9c8NTALC5ite/a8wrtlfU96kZFPpJKQEduVFkOX1sne
NLuFqLy7YQIrerxODhEqP5/8c5jmylJV4NxC8izHGdvI1rH9bdYW02IwkaniyH5EaHpHRa0dvN4i
OluGJreyORlvgzc0PFdPA97L5TwpCTfSc0QkWCDTQp9XfouXwkoD8tCBaWBb4suaFlesCXQO9e+O
8Mx/KZxSzbByvlQQt00tEp2k67O4GXsvSmh4tds6CP8cKSbhAd0/kqSmyDJea9hCOjK/xFm7qSdZ
fVpjMEI/0E3yXlN3bKo3ZhTJ+A+RS9kTOm+KeKHIpuXYc0tH6ntDb8+DQ9Pf7XqLjUXiFqza+u6i
/BE37KoDisEgPsJivqhLWaFuz6O5byGDSxg7RmnbcSvczrqxTymedMrYK5l7TSjNX1CfSaebwPy4
g6hD48oI+yIjCnNb2NQxUYTVsxYeeFTg5MSQUlVFTrNYWNkUcPNrPvAB2+gVFwImexBXroP22dBq
HT7rIXBZNnrIcqt+Xejs3t/JcaT0DHd6Y6gEUMW4d0HiuU39LeFTBqWNALDpcD/oHJTlAxxY3w1y
kvzEAOGKtvmiKNpG+Azt0omiMpCICv0DlZJQ/JZ+S5KxlVMuXZbiY0VGroRoT/8iXrmfye8IK8eP
54t168HlX9BphxdgMdTHg88fzzhzjzDpnPKNAzE7VEkqxSHL/E8t8zuY/pPtOLRSxpdzJJwb+WII
3uJan+egoTaPMdeI/UdTyRzCJKUz0eITZ0iHPMLFNhPyDLPV9HArPM/FkC+ch9TdfTtZAhmq2Ke5
FTD/V5rx36bvIH9qTKBlt4iCk3KX/BqhLm+sE91cHGi7OTVIe6b8yh9hIgRjqGbOC4lj23JGzQs5
P/zP60gAZEzqZ4skQm6JhB6VOMrJiEwisjVHb73fPZerMnQmuyberolR0Id09YjvfyoGzkHu2+A4
priiPgC7z/usdJenO0aKjBjoKtJrYWCVwCzHgHrg2/0+1mj1YtqyQJ3kMXtSC8c1XjCQL0+x2MsR
HCOg899OekRH+Iw+pKfhCi0gY11JFcZ5MrZuZuK3RVKdD2brwsWczMw8qHVtCanip/yvSaDMK+xD
iVUjuJ93Iilu8hsqe5h2uZMl6qxihgYAUG7O8V1DZAI2DQ78yQGobn6zRe64eoQ9iQon566rKGML
Sskx/ovWBuBCD8jGPZwKekGuW6QQIgV1GpPpOdlSlQZ7B6lUnGv0r69/uA+3ZsH2U/zJhI7c3aiP
Pvmnv7bOcVOBFulBIld3h/CsppIXN3JpbUDCu1R97MlPFZTsRC5grT1bDCAl/WGW48rDeZYqFAMu
dv0mgkjue2Jjxlf+3FhpT8ovCFn0+vCNHmyNbMemHryGi+f8NDj2zIF9mmSRv9ScMa1R3Lg4HbqS
HDPUKTKd7o9MelABPzJ0+ruQKYJiAc0+T/N1cr/298OgVU7Xe8NxIKRfxZ2rdlVD+JadiJp/9JPr
igyQzWlKWoiCBGsZ7E9AwBVR6Y+cNJmdmSrwxn9yVVTxK8IKXxSZgTdcTmvhPcF5LI1DtwtyxO8N
W9wSu63mIFC50agMdW27NGl7i1dDm7aqHkeKa2l1CcL+vgMvz6It4TwZVUfLxMlEohJ92qaD8tQu
yHVUiGjgYk9dJ/DqoP5Mc1ysQH7DWuDEuH4BEqCl2LNVCxAUsriDJlUGlezVs7bipdkoEcdZcMSx
+xGJIg/nQo+Mpln4XCcJ9caxzw/uN/2wz6vXvsCt+N76Ajb7Mj6cJ46mvMKeSJtyzdeU3krDeV+c
vVDMRYQdVTp7gmBGkGFOeG/CeexI3mCiJ2zW2xZUczlsWiEHd0HGVZahILOwmiJS2WHm0Yh5/uPl
dkoalHVVA/gya4s3UvJrtYt1JT52PKZL3uqugi0u+LkXBu/yBSj/JqvpYmtvy1z5esN8xru3L7Dz
y4BsRT5YoeqmNeaJxKx5XDTNKfJ6Q+8neqq2deVAlnasWlXmFbYn0iqKSczztXSi2f/1PgB/PjAF
uZomQvKz8AQOCT6zo5Eb3XJ5B8k/LnwcTtWHZ32LDo16RVXZOps+PkxBLSYN5/Cq3D1yLpwsGj6Z
ft5uDlcl+Aqo+KcJbCIGkO+KGt67gIY5vPgWZhn01vh0Aza4KiLQ/D9bwY3FNyMCisW9QwhJkAey
PPKbiQNkxyh9e92bGWS60VuocSGOsiJLR2AY6I64s31dt6IHri7vzPNgwKXkN4zwi5YmrYJvjRcz
sGcrUDJthxHwiZ4BVOXqxYvCheSbpj3EdCUbSykLLGY1/++z5lXC/ej9cYwvIJ+Rnad5qWuOVxVw
BJTsfNpYmXN3JDW5j7orGTrrlx1DDupyARENGrdzAZOa2w2V5hsKYVlI9vveOBifktmuFf4GMSq2
KmE1iBMG+BMoRA9OgTSZaoz4CeP0BTNhnINqL1Xx1bNPYyaCDw99YwpsCLrjXVXpsDHbTL/25/g/
9J5ioMhxq5xWfxon7GSXYUjsLsXK97OyecJ7Vxy5UPZ19A1AoOk14sGJx+tk5FJBSi1ts36W0gRR
oXYlveX8TvzfcmOfcDNa0V5Ou5Unx7UaImA9LLKvhgX2kMbIyTLOdoFEfPBGe+gsA7ZwC451ZXE1
bks6F/MDBauuHH+Ovcj6G0LfMI75c/oCLELVnnIJhQ+yO9dqIAZMeznG6JYKZa2YYq7CZX4pl9qo
hFQMypNMmajOIZsibxlaKjnJVXPqXZN8XOjPLU1GrmziZ7GqF+87FSLB5CnTuzrgVnaiSGV3uZYj
9T1C9R5xDiAopTFoF/D9k66Px6Ky0e460+cWCdAYsifa8nkH2DZpmsnGVyntpm8GZ5dD0HLKambn
f4SdugUfOd82DIAUtrk60HlrLtaCFC5wwP9WqCymL+gYsRD4SytUjyvc1B/pW1Psk+rZ1IAdtjHX
Gx89ZIWyHpvQ9K9l/mwX8F9N+9zoc9yik2XOUtDnDxji705mdRf0xc6zUgRCe6W6cyLzBg4i4OOL
6iqy/egq8kZzTQDGa9YR5WihC9Pb/g8n3lq//YQ7V6XUqrUyHNEAQe+r76Ahmo/7ePHfMb6l11/s
en5XY0z1js//va1VkH4TZFScOXvZ9MnrGoBi5T0o7SLsyGz0l5PhbDZQASUjI6NlW5BOwfJF0ScK
g+pQyVnMixmiz+8HPtLMkoMyU/4rFAKvC8pNUhUegCQzm1NTpdSq7+J6YWmfaOmgGFP2bXEHN1SN
AQvpARUtqvnk6wPatE2GhaZwVakJ4RQn+X75Pcjqn+trd0bIaSQaPHEFWJvro9xNc9L07sCwk5nH
caSEjeyxsOQ123/wCzf/HOy5RB3LuaZ2rO0MImCuYTytpfs6mQ6Vb4eoTAN+s9s+sOk6fFTV3/qT
0636WwuHvXv33aFOAybzzF9ydvurFq7HfjemG3BO4Bah2vYm3uMRc57b+FlhG8ErTbH6zSVZsBD9
0qS6i/zLjHC/Z1nvQsa3bPnJCBAZxos5ScV98TSnN7XY9lzcREwUuQ4q9e7LQFkzD5OhPbST0VpA
C2+/qDE5pn9P6FY4Gu/OJ8dUbMdtrx8w1GYQlwx9Z+TohIbeEqiSLBKcxv2zXBSrkMn+EEWHMCFk
LWB3nzhmJOTF8ZfKGzUTMGBmOm3v6Tmc1T3pGaQRky9P4cp8O/m1PloP997Oe9IhAAfDpTw5/jgf
7mw7JjdzKr/gcOsxInr3rgBBYwTzmMo9jfYwa3SQYBYj3jXYA5QLYvqw73DhVwWdgOt8DkkHctmF
bAV1nXJj0jH6EaVitpdPXZhpqW5HpiX484hTRUOK99v3IekZaCA8fH/Sdax8YkIxSUo/7BRtaSUy
WxdoKS+7eNqKawf2Eycu+zJuu8ZGLAuN+UciEwaMbHnU52wUSTx05zAhzNQ2wzc3ndH0L3jqtHAO
QfzOhTOCa7mytecjB91MlV2Q63t4AsfYiwD3JmwZ+cE4B0xit+BbJ/UnbWTsJVh9pLVwpV/+PeIF
Jo3U2FGh+T8iGev9Nsb46vNDccpgXTa1jedlfw/hvAQtPSJWZzJNiKncJI3wyjcFyNX2/aZdcEUc
ixieCDQTXSDPCqM+GwWd1NcCJg5cnkQ/SHnxndOG3UyeSXEVRUwjBuf3qCchdONo/Ve3+hAhjc0s
6UXuSDbV6zuXKUoz29KJgel99TWrkBJbQRD9Hmt3B9zuSQ4AYy80fJKKNdCIGwMC+kc1+ImdrBsf
j1kEQS5vpf9rc6mYDc2OOWgCuMq6n63IH1qZ0YHL3unAddJ9UYMGvI0sYCSbq9394YPJSY3pVXQx
/IYoM2jnaLkCeIXpxn+Ov5Q1mIC4YYIDQENZ30pXX/LupkSqg5mjuuTxuHLI/LX/nZ75ojOtt4c1
AD/WKIXtiHEVxfHLSYwrfhzURnmt5N8aWM4RTsR9+qpzCV2tNUWmnt5JoWy7OZ9KtEok7tiGD4eq
y1/ZBV+dv266zQK4Mc0YW9n6eZJ7gZ8gXuzc3iHg5KmAPGfC9uqUrVlvgXfvI6oYiSC7kY6CckJT
oDsT08jYlqqronTecz8mtaj8+Avd7whPzuHbgLxAFh5KUWmeFoyGhXQnGePqzb+Rr8luARhOtjfL
hhF3hugskgU9zciOU096z5VB6u6WdC6zh3fhAKqR1BJeu7JO/vbe0sQK/hvfj1QUoSll+QvtDq0V
DKgJeHjP8HJRtIi4c/KDDqVY68ic9ROhRXeBm2e6xZQzVdNv3CaoFTsGjBuXjPHqdAa5rL3Bhlql
F3PhMqR7jZjT/FPgDK1Zt3axZRagCqMrB7veQ+xRU00Dug5YHXHqchHDWjthFw+mh0talsNu6sjR
k/pCtPn/WhvIWfxSBeG9u5u7ZEMO7VWRkiRXlH6MR6MH/mhHpUwbfYARE96NNj5zhwHKqeFCa19S
CpjuTIAqPfWYUefp6WNWdB6R/Q6W90ZvVKF2w+D2NSwHIAeqX2ph/jwlByd7i4Tbr/gPU0Y9bDwi
kd1/Nyg8vAKEIE4EYOKMJJ26vuqRtWhvyTmFo5rvX+jhVFV7vbiXQghM7OPjnPNIqIIv21IOKx4w
JYiJgnAmyQuv+/LzHQsZskJ3yC8KyoSA4o+//CR7ZJE+zKbaNPCc6RzM/ElbENrnrt/AfcDED9JV
2ehR30NaZKYHmerD0XRCAV3cNYz7wercAB66YaPWfP1MQYoarIYhlNgPb1gfr6DtaHSXO7HS4nBe
i8vF+Rlofu2Px0h/9WieXVaf9+yIIqjUVtWEl7qdiaAKey/IJK1MO0NTH5Y7DlDKPTneUi6ZK/vj
wtNDnoMOyKigdA2MZMwge8fn581fLnoh0AADMCCizC0Gs4aa/BKBDRobp/E6WytfkWX8tRwuhXqH
8dgNWqb9LM1YKXo0m/XUdYTMvTOwibzwUDrctkUpP/O5gNmiiBEzFPgHbVPoO6ZtxCoY2aOLPTMO
9MPqy2kphlkROPfjcEW2072o8blpohHumETelfSMAktlIe7WnMr6UBanQzfPx+mwOdbdVbqJDtim
vK7B0k4tU3FcHhWo6nrB9T8Duii9histxYAGC/rj6QTFTZLXFBx3kDy0U67o/NYNiMYsB+n2dIHZ
MU3Yykc1uUpZCHipmBwE5oQFyHtcRClA5tpG6G+5YLCPs+li5VgpI1iuFRisvhwoeK75baCwx9L/
b/qp7DbABT/8nDjucJQ0FJ/Ao4iXTrxrdi6QbC1K4wi8Ic0BWpIa0H7rTSTyK3Gd+/HgGbbkuQse
y9ltPUryxTedFIj53ilTPYJcZap5pQwAvU+SRfzPkMWUes6uRzqLMVDBTNgSuwIQykTBpE01br5e
IM6WCv1TvWTgO+NA0d0r4zboX465DqULS33yCjCZFPGGozKlDsoaS2ExZWaJUEvkXXG/cHHiF6n7
YJQTYLb4iwTYmuuosvtmDQ2/u2sA9xm50E/GHPTRg6V6bavb2Za0gsVQ+DF4supvsDX8or3urbSE
xq8z5wC3faSXXyRMiPs1Ie5WefKDG3U9p3Eou0DWXfE8aHYcslDUmrr6ZTdl4GaaK0kReX0Y82ur
XqfiFyR0ZrUUoi0NNtR2XX5IMI9jnMNRsa+NKVKnd26NbyXP4g5hl06urMmrLitrxOSLedadIY30
rhpRVDFGnCJfyGTpsHl7lIdYeVIzxE4/0re/dkQ/sAawcLkWyKL/WO53rCIDyDHGYXOjdpTm0Mpp
7FZ0E9pB1P7rcAgb+TjDErIUw0yQNk010y6sOvVRmBnNJ6mdVnG88YkM1jCUzGs2NxtKitIWNzBu
R58C+22ciM+VcIAWJEMgRw5h9oms2jGmO9o4Xs++W8M8Cif6EeILSjCqAtzmm5ZZm1sTBrVoi5Ua
35NyPnzllMkWKbOV5WbpS3ji6VwHlXKOcJ8gNSUQZ+KWzU4UqjRdodWsTzSq3KPcA9DpCkTt2GOI
YhQCXdpqU5lIlTR9fhD3ZrKnu3sq+jMcLjIIuPZKVgJ0fX//4Ycb3wG8ez6NGJQ3JN7i9nLrSF9Q
SrnkDvw32GkrxWqBKQ5twB0Mr2kFFX1MBlomZ00SbgAbQLkcmOXZ2ACtO7aqJdDMF7BSyHy6sYaQ
JsOwI87SYT727l/x+/PWFB+CcCGqAvG89RrKmFqbDAHZP01430P3WCH3CmwVS/OqGCpCrVBscEEb
haL3bCcD+WOyx+1Hkm/j6NTpRviXbunCUTQPxUSLQ9o7hhgKVcd2jiY07IMSlOAMDgVo5NoigwkM
t6Aino+pwp+DdJULod0Q+u9nV7q9KN3WdgT2N2BPs81/FnMGA9WEoa07zLVEWX2ohX5dBHX1WaID
0Log2u0NUoEKmGMACvlHvIHxOuSaMoOA/8R0R23UDnlDxckC88WjI35bDC2dXH/GG9VCb4/kvpaU
NNnY5gPAMR4TNUyLAML1p+zHerXm+T3c56wscCV7QFcuRSlp+gW9aGUx2yo8FnMCkk3lstFgXJUA
2oY5kVwILR2DgTL/jJjmPWStPp633Lx+oQvMvb/0YZRv8LQSNr/MlUV5IUTu1n7L/WzHhXA2Lag6
4YXW/ocsEIjCCVYicFSJWDxxUhpbGRYM78m/hv9mkNyhSdc/kQRXCK6SwutPVCiCfda2LTsxIdPD
nIh9Gw5H4ZFXCJGBKHHew2fL1/sm/IxSwXQ3faBiLLjQp4SBud+hkqilk1od/0oKEmSb8Wpq7ox+
h67o2iI1UzVUEb/yrHNH8PoO/78IEc+ertOgwZ2WIsWQsgLUX2Y6shknq/bPk35pxKgzddMEBsbZ
odqQdRtxWZD/h5Zvd+V1sLSbOss6gC4AY617rtcnD3a7fUv8lUSCK4FANny7kdNZzyAFFlv9bcMP
IhO1g6l0U3x8fLTNFU+DrvIYpIQvhKqzNeMIXDSDnaIzowfK373iEZqVsnd4hIYaDeOfQvMM/Vkz
dvU3ADkMiH0Yid1b6KzQmbOSq1iMzhIYxadsqj4NwnO0FeIxYssvXBPtKLq0QePGUSzlPLL+M3UN
Ri7Teju5PG2hOgSf6400aejzkG/ichqgvbK8yR4G8vN2+ryb+POwNB9Ph9lCtE8gp1Q0KxTftpbB
3Y8jO4NctWNlVQIijHxgBJHMgiTk6ZilpegHilmAB+nEwpktD6mHCBtSNq2WSMiBHNnYGFj0iHal
RZuV+d4rk6UGHCnrqBB0mvZogTh7gcE67yUVY+xV52yyDP1fEUCfNa/KTbipa4LW/kP+cKPWVlXJ
n7nIopRLDF3252cPn24maPmHk9z9H6Wx/lO03udDOJWzq5BmC5p10MlWWCwGKivPjaeNS44kminH
z4APvissx1l9qDX3gLGYenkJVUzrBSMnRlQPrcIqPZr9ikR3ln9/VJpa7H7dcgjzbQ2VjDXRIkDl
bSeKr6EcQlsPpTynRZB6jjRcWWyzD/KwkG1RyL384qjDxDW6aO1ndgTZv3BchUrsYTTUHuaEeVAV
zoiUQuPayUdcNiRVXhjGvKuP7RnGWQune+5A+uRgZZ7mQlhxicNhTyJz+IVA46w9Xxdb2mxB5knL
XUnv7/IxajhATQugk8wIKtQSw6bP32Flk7hntD9G4yyL3R7E+4SJgTRImw2vQkMqzK+zGKjvv9FI
JJo06MrbmIOcAGH754Fg8SMt5n8A4n5JZaKjgyCxCiyMStI6P5nOaO9TrkmQVFUI4k+3cyJrLvFa
6Hr5HgYj7gyDJPMBzkIqUpJysd19KamBkqdqZamqaruNDNe/XaJV5JDZij5wjgO9u072QzXFGMtG
H0YJGdo1woj/7QouRnEHCvi//LxYUxK8Nl5cfxM2NsvvuFohrumGYW9/AhOV9P1XSaap/cnXBc2/
wYNzIT+8tGyZOBPXlnwzGjHfXejFetLPBg69xJB8Qt7Js4+j2Mtn9FzHSCfxwe93so2VvIwR2EPI
GIJsW5IJGANDmivAo6oiVN9UQmFJiDtuPnqAp934KbNiyPkOVAoRiKP5EZQ3y4pQPZJRlO0MD87N
fDKGdcPh/qLZF1I4j+JFjKznbhgquGx2yJKn2p19EE84KAfbKaMx3+d5bNPgeSI6fSnInVbxB/rY
MqprwSpMnJEj1xeFwVYGc7u1i9AqmPxFb2SFsHj458aUkvqb+tu0Af0eBfSzJdwVJXPz4HO45YLl
RyFUiOGlsm4pHnPlwN19NXfLoH+tRew7RemqMbAS2pNidAvugRJvrLRTQbNVFpJq9JINhUSXd2C5
`protect end_protected
