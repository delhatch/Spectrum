��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����ս�Mm#�&G��BaUG����5R�ۖ��Xyc��N��2Wv5�n�[��|å�6糕�=d�����Q+��4��JiVE4I"6ya�@�Fwɮ�V�Nhݽ���5Oߍce#�)�<o�]��ͬ���T���P���W7�}��{������[����qG�*9C��~٧���ͮ��|O��:��)~ �ʽ2�+�Wȿ��� ��;/C�����K�}QQ-�8
H:�^�p�
�s+̼F���2�9���}lb|���|��$�\lq��q�ɽ)�6���1;2���kG~z(��:���9��~��`�
��	����>-�����~����������Q{&�4��qʮ�{#��
�y�C��D��H柳�������箙�0��\���C�W��Ǖ\,��\`SRt���n@�T<q�Q��^��n���i���`ߙ��q03<��i^*�){����Ҡ��}�
�I#��㺮Nk;y��]�i�m����}��gS;��L�y���?s�(2�lx撛<�t�`_�w����G=�;э�M�e��:��C�3�d��sT���F��~%`��cI�7C4NL�6�a_�����/���I�`塚�nߐ0��$1>��9D��mP�ّ�R����ة��a�{���ȼ�d������x�uJ=e�Y�iP�������Uم�rb�P�O]�$)��I5���aR��!�e�_a\�8'Ή̠��6%!��(K��#�7�ڠ,wp`�Ók^3}���E�DO��{ࡾ��C��	���
��wK�ơ�>����X�k���,�܎0��)���갠d�5�j�0�� �d����8�-�����'4�ҹ"W��񾭕@A�ʤ��jN2�n��v\�}[7I56��~��l(S'�������OU38�����$��n������	0��i�~�R|�ь��P���)7*W�p}-���tGnK5����$6��n�֏�Y��M�l2��D�{@����h�.JWn$�7��ٹ�a��y$y0Kԝs�Nn-~����Y��q�W�n2�+�RȮ�d���/�}D̖F�a�bh�������G��������W�
�^���s��5�)���{Y���Wh�N�d�����Uc^T��b�����V�����$��06��I}2˭�Ԓ�g}��k!�h��A�m|���ֿ�H���,�?Y���o������d��s���}���_IS}��۞�?�X���D�Pjn#��&����������ЕB���7�-j��K/���4���PО�;o Fp��l����B�z��w��|;����ag���N}��u������,�y&����;z��M���nQa�!�'iN#�7�������B�2�ɍ�Q������+mk�������,�X\Y�xg���_��;�����}Mp�|lB��
y�E��ʸ}J��AĀ���d�/�Q�~R����]�崔�ZPl['��w���E/��}���f����;�����)��v�r��p�*d%x�ce2���S�ih�����sUe�<���`�"�ӊ؅���|iz�5_Pb:i�уq-K�/Wp�������L�8:�g�I�Rk�!��L;����K�!��}��	������m�ZL�Au�Cb>#lN�*���yE޻�����ը>Kg���a]��I͙��Aj���6�K��8⎱!t7��-�����vG"�Q'��WU�y��%�H$�0���0#mjߘ�`�OUD�'��a��XقAr=�)g��2���ڔ0��dd->w�GH6�n��G��o�Y� �V��a|�}��o�n9,�6�Θ&���p)�Et"�/} �aܔd�K�O1��xpP�y��p��' �$��hLp��5pL���q����j���s��A��P�ol9��l����WN@�g�PSWd������/�9Y�H��9O��q����R�"�	`/��Z �&q����$w*����d�#�D�`�u�2R�1�G1B�V4���r�ffޔ��E6�EZ܈ԕX�r���:�|���l�ȕ5�s��eY�~���'��~~z̿�V�4e��CF�"*�!F��{����@Uv�wt�ي�;n�jF��X����=�@�$�>"��M<�em���o���e,�P�_#�U�ѫ��E�pPA,�8���P-K��9�CѨ�?y�2�Q6H����>%�<}� �@�]9�T؍�/�R�Hx�Mܑ9zw~��LP'�x�xt2.
f<�@k�qe��c�4���n)�)nѧ
©���Ϡ��4G���LMJ8��'/@����p��dSR�Z�G�R��bKuv� .�Qu�R(��/P0}U������)�4#aV����(��r}��L�.r��ڴB�PɊͪ'ۗU	Xf�R��}��4�}v)jd:;�I0_��`(~
��$��C��1�Ȣ��::��R�"�3��պ|�$�^����48'�����X;-� %���j��4�1�^=L��-�m�r�P�,q�=@��[kT���F2���"=y-1��[�|�.%!���jp4J�^|�H�s���^j����D@��$��>P��PR�D�����r��ͬ�N!ޟȸVdZoM�0���O}=������aV�St��]��v/T�Z��rF�2�x��.D��oT)M9ʍ�'����ݝ��5��]�)<��,N��^�u|�Ď ��c��x�arc"��K� ��'r�PH�51f>:� ��q�15De!��K$N�X��_9���]�&N�%�A���o�N`����I�]���K��l�)R��_����bs���cM9i� =��9)����n�tH
kz#YO��r�z��݇���6�N��f?���4@�o�����-h1hk��&��:�r6[��0���_���W���a}m���m�Ͱ�B���gp(�>�D��M�D�C![d�@����#=� �*e-�J4ȇz8��Yy+�S��<���B{7��n=�6>Z��N��� ��O�~<;X%Ҹ}̤���x�K-���>�����}��9��:4�&{�\G=�Ǉ��g�S?SX{�Q�!��n��t�,��E�Kl[#H@*:^�v-�݇��h�2B>Kǽ0���<5^@�A���j�mNwq]�|øR{������D�Cp��B
ι���Su�d|��Rn�V��*Vt�o"���hHgOaԴ-�8`ϑ|^�o\�/���� m"%�'Φ$b����=�9��_�y���RW�b�9Q�6 �ZP|CdM��%�����,�;��Ѷ&5L��Nq�������Y5+��Ux��TpqG|�:���#;0��]O��x�S�y+u�(���Ю?{z� ��]��z�8m�h�	�M0�+)�#��"hu�R��g�^3���l�(�O%]�N�P����o҂�ow{��~��i�_pVE��)�p;�`�L�@�c�0�S��]�"�K1������Ie�I灢����E�f7��D@�kY�M��f�cV6���Cj���p�Cmp�س/m���ĕ�y�pW	�i�0ߺ��������!�pa�vu�]��4��i��'���D�q[�_��wt2�'�3_&��/��ԈE⧳����5!�-�ga*�'��� +�4��<,WaU�6qiC��#�,�ztd�;���&����T�s�AX'8^�
�zZv��옓z�91D�d�V5��y�HI=}(���e����􂅀;��`�?T���ȴ�4g���\ �W7G!��p#������������Xi�~�M��f��}�2��X�D����n%�d�8�Lr�[�.D��i�֪�q��ò�m����f��{�e�x�B&MN��m��@�y�t�5�܂<�`��~��1Gzu�9�Ί¯����������yp�#UhmwU��&KI�~q-�lo�,���	�O[�
����éC��v���l��8��R]�݄0,���18f-1xu�
rξ�N��G^C��ᾰ�a\\F���y��1M5ς,���.�	ȠO�5)�&�6H����
��0�Mk%kX|)#�(�qnN_��U:�@��^i*��mW����2e�9p0�*kd$���*�½��w:ly�k�9^�@h���1쓕^���\�P���'�1�z��|�_`�dP��_椅��I��K�=lk�x�����L���& ���,�e;$�h�\�,����a%PD�¼�7�A?�6�8��ZP⼹���Vh�*cl��@�Fg[D����a�qȧ'���+�1_HZ�}��ثɅ(�#p�gM\�8v5!]���mAL,�ζ�dԔU���\���J�z#p@���<ԓ�|�Xy�l4��;���YeOб1���i�����=h���yX�
�S�=�e�O���3XN5�3�̂�Ly�-7sĲJ��@�C��Ե�[#,[��	l��B3�E�/z�8�����;��͚w�������YS]#�Wh����x�R\��>W�<�k�5R�̮m:n�F�4����G�g9�UU	$w��p(�P��o��c����H��E��o�);���ꗻ�J~Z��ߡ
(0���ٴ��(�#����{�����T��=>�����L=I��_>�Uja�k�~#LW-[��~�R �����>��o�C��N\U�nD���3�ߜ�>lN�A�OM��Wi�)0mҸ5�����=LR��@���+>����`s{�y*3�0�@5E�Y�?v�̞�r�|���Uz#�>�ezw�R�@	���u-r��Fq�ayLTL��J�w��Q/]��	�ؿ[sj�����Qn���Q���h]bw43��)<��V�1p��l���W���ؕ���r���+�����*
_�����R����������GK��ӱ-�gC[�.�#�����y�O��x���!P��A���8�%���e�� ���!�<��$�T�b�jԫ�`GRZ��.TJԩO��gJ�6V}�s����}�Im��<�``_�G��#���36T��41"�<Rx����}Ⱥ%�L?���6�t�E��'D�i���g*�{��	Ov	`o��K�1͙lw�*;�'��Lʀ�_�0�U4DՁ�=����lXV>���h��ϥ՚�u�桼���`�Z��D=3��@o�d%�Hm�b�`��:�:�b:�kV����&Y�
b]r6�/@�����p�W'}���d�+X@�|LW�gOf�J:�P�Z���hT���L�)��X0W��MP,L׃�$���j��	�L����j�����@=����
 �!�~VeILٰ4�]Rh�&�.K��Y�
�W��;���L�ޚZ݉W�݅�R���%�����A1�������ƫu�֕9�[�yf�~��,��cp� ����'O\�Q�(�[%4�$���ǵ�a\y����|7�+�AƷ���� �H]Ϛ>�⎱Ժ�?$�,2o��Ta�px��=@� �ۥ��"�� ]�;�u�M�K!�5Dp�&�S����KY1��sK�����$���;_�tg�e�<չ���{������q�����5cal*�$��7B������$���j��ˌ�bX�����#��w�XV���An��1�"�����qu���|V(]�#��4��>ߗ\�=Fⓚ���(XfC)	V�cqct�8�l+ESV�[|/1H$g��EB@ ;�ٻ�A�u��*�x�ucF��hʭɚ��ch���\�3%)*V4]�~r
> �hF3Y8�l0��G��X��p���w�_UJ���v	�A�g�uh�)]bu?)C��A���!����,���Op��s�fv#MsڎV0����ϑ[��EI�8M��6Vg>Mɭ���4d8dFtM[���k\l�+t�:��� 5����ɚi�^Y�����aš�Y:���Sf�"��VX�-=��D��z8�j),ISA��&0֊�㲜v�I�I5
{�H���zO�j5���d���M|��cy��Vq����xJ�wF��B*1��� �)�i6���%O�q����x�VN�����eI��Ѻ���+������"�	��U^�EŹ\0�o ��q���'e�j��,�E�5��f�Bw�!� �0�c������24��8&�+��k��ڞ�:�ͥM�����?ȉ�f�LQR
M��q	�Eȷ����u;�!c�s�/U7�3~r����M�a�����	K����>��U:�x��%B��V����8�!vR/;.����o��BW�z�L]x�tb_ V���)U���ß��O�]���kJ���ɖo�y�x�oKP2A^,5����,�D����{d����w݂���B�<O�&$.-������ٴR�ᙼ�6/<���Z�Z�9��M�Z~��4���B��e���_����ce̋C ���u��i���8bZo��$��XP���Բ�@Af!��;���ї��W�����*:�3���!{7NI۲qǤ�v��z�x«N��_!�`�X}���k��p�Z{u��	@x=f?��H��Zf%C��h��(ݭ�'?�&�'�k�)�%�U(suԮ����8$�l�_�,��U��m�rm6��	����>γe���zʫq�!�7  ćM�v�]�����������{�ؑ�/`��,h�udv�����}�/e���FbC�b����C's�����~�L&,-~Jq}Cn�>B��)��~�͆�?��HkF(�R�����T�,��cѠa���`2����#�Yx���rHQTƕ��w��+7��\���/�z���:�-�vmq�kFf)��q��߲l�ea����|�@
$� �~�:}X�w�K0T2��n�N�ۖ�l,�d�Z��7ڲц	C6��-�֮id�ܺY�j���>�׵!@^c��6�5��O*
wl��sbXr�vm�,�7A�Ѫi�>ho��NqiLI8��+�E�2����t��Qõ�!����r��x�Ϲ�������HU�>���H�+{{�t��(xmr�jӞ$� ��ӑ���!��3��>��K��A���C�ut�a$�$F��Ry�h�R�;ʁোȪ5���d�A*�W�uOZ]����U�P׭���F}"D��pl���}��H �%���6��|��l��޵8��#0�gi�	�%Ѝ�n���4���!�f���8���e�5(�{�I���U��.���5��O/Ĝ�.#3���$��Ɨ��d�h�����M��q/ދ�N �6�t	Ƣw��HaϽ�E� &qx��"�>����8BдԅRQ��� �w�K:�DӸ7�	���D*�Ș�#�G���r-x{�-����C�|d.% �v�U�V�4<��*�*�Q�ɰ�%�-ӂ�%��⩔}�E���JZ�Ҩt�P�]Y�;@�4��eJ�ȥ�\�B��O����t�!������-		�.���<C��\�$��`|���2Ln�/��l����L��7N���:<' u�S��	�A�B8�]/	����<�9:E�8-�;�M�H.��g�Χ}��rI�}
��_yxE���;] T����]pr~����F���u���x{v�k�6���OuB�פ:&麊��P�w@;m�������5�j�� ��
�QС�����k=�����i�ܨTA�o��ܡ��^�3�A����)�8ƪ�L���PP��zq�p��A��ი8�В��NORS�� p�\�f���gR��Kq`V��}�Y��wO���8\"%��խ����^[
R|G�xG�x�#�f�8�T�Ó��r����x���a��@��K��Pd��F�=�SXG�]K<@�r��V۾�����gᴁ���k��&�*b��>I���C)��3�+д�������O�g0��+�甪p�.XoE=��h8ӬJw#��Bk�k�:4��F�r�j�ؒU;�L=���MR���fC���U�|�n97LE$��2��kp�����EB�R����6�u��� �����m�)�2��b���Γ�ua�7���
Nd������H��7ZQx,*D�!/w�#�<UYdF�5[{��6"�j�WR��>8y�*a�޾��Z������e��A���˯*��=eB+b�!��%%������A�z}�g:{-��zk�L!�T��V���4zw�S6�\��Iď$1�n�~0��`N�<;�1oH�xA�,����N���a7�-��܉ox�UD`��_�G�)���w�%���2>��u�-�2VwPW���/�N8�^fL7�[A���� �9F�cSG^��=k=��Z� />�T�H��S򻪋�yם|�Rži�1p��L��S�C=PZ��!����#zI�iH}���;(��Q�+�����k%��H�L�I��/���*�����'D..7`�a:��B$�^1��*�\����qV �j�n��g�9��� vw�-��њ���-%��uD&�?bA�˴���9�<�f�e�*{C�\"�~_���Y]&�@{�Z\��tJ��	
�+�L����C#����Ɯ��a�o�37=f�t�m�����vF�O�P�W=���Ń���*���cV���m�S��K6����k�Y�/RvY���ˋ�M�j'�gz�P��H�Pd��W���'�B�}.oy�fwҏ�S�$i=�/�
��Ơ�r��n�R^<f?�Y&Y��	E�!�R�R� ��|�F��OliH��&�����	C�aa�Ս��[{;b;D�WT��M��4s�N�d@�/w���6�8�8~V4ۦG:�"�)�����!�D>C�r#��}�3O�]Nx9�Ȉ���JU���iA��ċ����XpT'�<�k�޶lG
{����;���k�e�y���f5y2@�������g\������˾�j�@]���C�y6���-�c��N��&I���W�g{=X(�o��!���nxn�l��J�+��G�&��"[�sQ�2�ab�O�w�R��췱K���V�1��u_���vy��W���w�褁%*�M̜�H�X�9.��
I��t�Ȕvf�&��&�]���J�2�<�b�zn��J�,�Ӝ��>�F)��. �rP��P	��?��.[dCǜ�Ag?��T�잁qF{�	&��q~ŶQ~�cn�N�tJ����z�jW]jbS=�K4��w��-�4h�8��v\�R��n�{a��ۓ���e6���}1F����j�j�ń�:iY. ԁZI�:��{�y���������t)7ǚ�5�կ1:t^lo���8i�%��������'֫Dk�����{���	@ʃ4&�%V����3���;��EyҶ�aٜtԧ}��9�[�1���8��aI�"ZUG��O!F�rK��|�2;��̒�ڷ��l$h78���v�]mU�7���8)��~�=�:6�`۝��ǂ�W������c!.�!픱`��Np���@��)�w��G1<${�.�:x �<�l��l�$~OB���E1���0�O�'���?WO�w��u]�Aw9�����8��N��Apc��^�����z��jԐ�r��iem�ŜT�̎i�<�]��¯ŵTiR].4����?�Ү�O��pm^��pJ�֪KOg�D���1���i_;�w��m����_H���
R;e���?[0ٯ]�y�AB֊���d��ѓ���:��)v�&c�y0� ��.�M*�S�M��ٴ8Z�kN���=�&(�����)=�=X
�s|�zƓ����S�V{ܥ_L$��r�xv���	*ćAS��JJ�"n5u�V	���wx��g��鱛4�7�