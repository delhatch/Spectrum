-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZoobscgJUcaHiCoJBpMA0LUALFkkgUfximvBBLlFKgbSEkUK8cLvSq11GArDwa7DYdDUJSalKRyx
4AAe1YMQBKMCY4KTZgEyKnPoMiNLhhN/bsJdvCpPc2J6yyQ921R+89d2lIvl2LQqYwZWEZAgOe5M
nvKSCb7+rJQcDJ6Eg2rPiUIU3EslTvZ6spYbTMImBbBLtMnGIb1q6FRReCiDP5HnsQQ8JhSE0LnN
/Ums4/zLQ4lLtP2hj25C16f0ih5Yv1FQQijxmE12iU4J17XivyGM7UF+T2+RMsHrFiz51pVc/WWq
HeqnE0OYykqlV2gL2dXQDZSTVQy0npc7igxVMg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
Hz4pC+iQxewEN7tL9gJqtAlu1EMKH5qnedLWSrHknofbH8zquyDfY9AJL7KSjRU2VP4IZ7fOOqTK
OER/KmCxCvmWlhm/RG6oCq9IBHZ4dT7PwVSPy0hCHbndGCVuwoQl+ymwIKCNIf+up/XBx2ZpC9g5
VrMqcR8mU5bxkb7PMZ1e1i6qoU6SdCpbLl+JuH7kqKJpqNmx71jaEwcC6KZuw3aeR6r+iKtUDmJM
+tQhELx9URv9qvfycIcnCwIfao2UNLjgNLtATY03BMZcIMiJDYX2+LVs9sajT/XaW1Js+9hWvK9B
55BDHPtMQjxSVJcd6lx3Zq2xejFcvnEv5G7YA1QSlEEVRrR16E3/SuxDa0kMmqm0x9lGt/+0RlRa
8XpD58Q7OONWysITTrKdh+xIDU+ZOyNX5E+fphh3bVGDkr4PkK2YOYcGYQNSZwuFuBnx7iE5WSRD
4lO/8cUSMnZEIZZELOVakRcI80AHjxn7eGticUg3dHI0UUqxInNq7/myYyF9lzqIyoutezCyZsIt
rOM5XxzmV/3kGoaeH/tEVGxzH9kFsOTGNFD5uCa32RGRFmxT4PEzJuPkFw389TM9cG2NTGkG8+BP
Fmepi3d0G7bDpTBTAFAYyiQzo4pCSzjc/6DHXvNGKEnvZJAzNahKs1nXQANY8Wmai5CByyu6cs4A
PCL5828QcJovhco2y9eFiPVhVpqBc3xx8G3lqG6FCijIHEWmpAnPlWZSTtiLJ55wMw0Yzkb9m41g
BZ6wqrdNLFlU8hoEA6+ZRMBGN5yhGvVVD6uaZyuY+gawOBw5BRR2fSiSdl5EfY7Q0olv3oq5dFnw
1nPslBtGbX+HoGm2AxEfNcUe+vFNheVYx+6PFQkgBfy5Atc02z0HRMDXIzN3TtfHpusatizb3Hk8
C8TezAGa13shXqQqq/TNK9yHT7CtHopVvp4dp3itSBTq35V840MGp27d6UbveV1fbccfZjwb9bzR
P4l3FUUNje7wnmrZSrSqbG+0rRVRj6pXKA4XefypRZUDS+LEBnfeOzPVPZNRKfyomqH5NgwH0Fg3
YrHnKKmrU+/1a1gvqm5sRrmd401hRaksoHhVhAAtLD4iDFfIcuSFCjHK4ykyX2Bo5m8p/z3G/B9o
qM4FC5mQYuneoRSPIuRwUlrA4ClrUWi++RnYRktSNGWeqoJPMk58TiOb1vVH9LGTsMIlYAugof/A
yuywNEDt+3oT9lUFxiJs7rOY9kf5RE94MgZKvnhdmgBHuEppJuhdE6oItrT2n/42xNSMbG27X4N2
3uPNR/cfuOsiGL7TTW/Mhd8tTVK3ribWDk2rZygtzGAZPQaoTvUgKp96d9/XJ/3Ok3GJwvYDNyvD
W2BgMPSQJ4KgkhEbHzn8v5/Uzv0Xsk7cpwC9Yw8YeGR9Ip17BnRO1as9EFJN1r/qeaCzfXEf4lzk
rQZz6zcQlAAAv9yCi+mDk3zepwS0X0IFX1JXPw77YkwEb/jr+Vd/LrNzniseg6JO9T+E98GprCQg
w5NaRA71eLe9eVcJPp0WY+FN7H0RBEZfUIf+bbrbw5H3lpbDhcQCqSXjdL29EOcKbZXuSlxOnypF
EVyL/t7QDHAWplM2iKGfRx2dRKXPCQcNAeqI4g15iypdNvIqC2OIaG5Yoq5HFmsPsMT4tONWMeN5
WBqLHRu1dzNdPsGbKsuFnmS7g6fvoCyOFDi9QzxNLnE6XevBgO6D1h1ihJO0h6I7bidruyBf4Zq5
2EKTvOTGskTK+jnfJ05WSz3oIUTcSuuoq4aacUFxKzigi7K3YFhUaSRhh+dQMhSDetmbCwORra29
aSqLOrB/IrKEkXjMseXxPL9VS3YedwqzfforoZVnYa4guGwK6d7/SYmwOjQ0QwG+iz71h4aU8c+D
8/aecwVGzffiflM8jNs8k+wdjGdICJ+WU01KA2fjsej54YUoLgnGHF3o8RbyLRHQVDaIA9efgA8R
ufFsUBXHXTYDi4RFeunrcyswHp7smXDngs+FDVRN7FivEtQ2r58+Fs3IyKE+T2wrH4uVJE/KN+yA
XMm08XBIRVW6UMEyyNSbK7ZfX51UpTg+RFi0TSzcf5fOoXZDYOiWnHHtHyn+K+yu8oCjJ5fes6VS
sjGceQ0YymiF32pePhTQlAYIQkSpGNrSJ/WxeFD80KNSnsaMkDCqUw7v2KfQKMltY8/9nYFtNTfW
3zp+Na6euEK2zO046ABuGBtYBzW08iQ6NzqMGXLbGpXd4jfbWrZ+x/HDa1u49eHOHqgCc2mWPyVg
lT3n43vh1Hm9bYcfaQp+N+IqRawGDZ7BZffzI5BweGvu3VcEGhhzdjAsRgLNU+zLJg+pmwttew+m
sZH1pe6shDpLtAMAstk5u7ChgBkGW0XLQnoAyE7LnFqN740gH0xAEzTkNBIe8HYGzBSQsIopYzu0
aJnpdSDtyzGlDkqYFdy+oqGtqeX7u64aKI1k1fcDQK54wzEHYwL4VbJF1E906ck2dxlpOyTxp5mV
UOzLjVRCfPNuMepsl81AVaw5DPjjQ+FNHUgH8RftBToN1a7UhKWIhQBi4DpWSl1apl+dQs43HMD7
BlG9aMo4/l8si+VFUDRzaW3LPUfhPlxymbZ/vIDqu+Q10erCKKkKef4OPMRKn//1Tc3xTODczvl4
43ZrG/z5+0aYGX8YRIn8geLuSNrN2znmPo9uxyiVS9TWOhzWVMYHPpTcCbSCvpIbj/ZReh7TALTJ
DqP8Rawy5ns1ODo2nAxtv0MYOxf6CA6tPQnXAuKf+gfdpF0DSnkn0fuoplbTg+o0xFOUZNb/c87F
epiAK+69d5z2UJKJDbz53UVhkTCLUQqGDqd8y30bRxo+jagdpHkW/U7fkaY5HbNpGeliDAMnT5f9
46QdtNWVx7hetEVO153w2kE2ntdeSrB6Ddwx6lXPYbqzfFEcniUIL6H/G/8wLMfhz6Izkzl/q8T9
0EDmCqPJNTNRmWhgr2knfFm6vFSgabICd1SXJk/SHZFOBrLIJ7DuWhBeCZDaRy5gaSFcVir+XKIs
uShT3lTBU3k7SBMnvyXesMAYA8zWfYkJEhleDN5Z+wSUH87YKKSjvcALQkEjem7J/qHURoSip1S5
G4Fd+OGoc6mMbeBNap7ORLSA74qbot6m4Qh9tbvThOa172ZSZS7aKcOi7FETiNlD0CrSG0giyjQ3
0LzhkHpD9yI8tIk4wr75u8XXKxzxHG/CWgwZ/McxYU7mjPbzRHTSpfINX17rFBpMuad32VjkYOTd
77uKWV9Z/zmzWWqOzxvhwHs9/aVbHJy7acSUSPC6pIZT3CEO53qwb3fZydJCPgnO2bgu2LeFdO++
4r67v6ZypuIsFNayiVzI3TGr9wVnhthM/yyVQs/zbF3ubw+uVSNWF52Vapkk3MNzFOQG1YaZHOp1
9kaqB5dzeTytajLJdPqivSoRQI1zAWlND/8j0dE3z9ABwPenXVpsII+vOBD2djcxUrDKt1A/HhEn
bgHX7OWEFkwTsX1LxpFS/kXDeuc4Zh11bwY88qZt1qY8iOcNC+YKwPzbFA/4Lj+OZFVV59lkRzmC
qAHidoWQaNSSS2wUptfhNqMX25SfWZvsqzYQQvR5IoDf9MBnGJ2X9VeXZN4DuLLmq9t2V6eZTq5Q
C6bX0reEdKmA4g4nyd1pn4mpg+msdLmYdPPYVctqmFGFg/2+CItnu8aomlLKxHGRPo0OUklutvmG
XNTkGIZWOqeEcvF91U+kk6HOe+brSlAFkvBroGi+xTsuVQNFxwDhCHLL+qPTLzzJYeMAum300BxO
m4kPbgkyX6b2OJFzS2g+ku4t4rahYD3mjghIXyTG8mGoSFvuoOIXQ7XjrH37PUDVcsH1Zm1xK6vZ
G7YfXZu0+tJtUZGTCv+pElTEJ51nm+5vNbRS+LqTngVZnCXGTsgX6/Iv6q9OK0mLiPajfVuNqxqz
SAlC3ZChAYM+PtXy9RO7bZ5niptRsKIqqvctdOtVxgUBFyEiU9d8RZvsFp/2jiFSTg/v1B7A+Qak
iltMn9xie93ep2K7bWqSVuT4xNF89b2+eKgswIjWHGir+0Z1QK9VOTOvyZcwab2h7VS9dXl4XWYO
2KLhQEnx1YrRqyANV5XxtVBwVEnfePyAx8MBMkFbeHfHFDirQJhpxc6Us43B8cd/sV9UEQd1FsuT
4LF2qva866zS4eEsZG+ylb0w3seGoOvNeykOxzjmLpcsWrzTbkxVMiKBn86TDfOG/ebWoO6Vjgte
OcAamRCBelKERS1ecobDZlBgeSPL+nft7AE99Dw0oIy09XRxUuagH/zQOAJBmRsaFyIrnebRm30n
K1U5DQemqlQDOagDnc1NT8eA5AC/5kRlH1WHG9Nq8VE2BaMWbLgkEr6RXRTodqH0ya+/qJUSV65+
xatUvlZmCYuzvizsNsPpLjVfIvZIR+rg8yIuahxhe4ux/bVHEq2wRVgHkXMwqf3BX2sx9cR1iaih
eKlegAvJDbfVF4rCIGaRPocIPhqFvwdMrqsd3ei1SDuqfR/I1ez8heO3uPEuyc4V3t4eXVO0xZe5
gv0XfR+1eqS41FK7k+8eEVfgJvkQOD9VLky+s+RdKOr9ifwhZMF3ZwYf5p4o9zFeRTIR0D57M/zl
ZLghfGVfyzgYkfrvFSLAn/uwkvTHlP75Zftso6qzQdtlkDdmUaNeS35zQKhKk/GXJ0BIrwcgVr/F
4QQ5aF4NcbntOrsN36c361EBt9fFd5cuDb1mEmGEgW4y3D2tjYobi4Tj74JRcIS/+rCfw8NcDZSy
+QUf+vx8twgqTCUhLWcz+EbW+lfxOejrYzRzM6EKDjcWJI1qhK3XAC7ibVexvLtGSdPkHWAXZQPR
jeQl9aZyUVewsb+iN2aDsITkQue4HZSmYUMU8ZehtsUShdVH4/fNB/T1c+HjrcaEcO0orLTORHLr
NG2fwNvz+BaJqeRU70BBEh3P9eaAunR0wLKpziLaFI8Chu9l1gSZ/wOP0C+et6SnyTZk0Gn7rRmQ
vSzhpFXkhDF++wY3m9vQepgSjeXiioEWkgPS45ulUtYP4eSH1Z9sTCuotKj1EI18vqXnSKYZncF5
DVHAoLF64wy7M5cUc9xhrUybqS+WzTXUixwVCFmastfoqTRWeqxAJda41+CIyVmzZBi8FtQT+IW0
/Vpe7HnFcPy/dpTA6IUcnD5HgxAEo5BmqvgZGvPyuMRBuzkc7c4XMe7vTYCXJECVzTAAt8Nd692y
6yG/FzE3hpzuaaEG6+d5j6/LLOaeWfFERF2smc+rwbGxS4OMG3uBSTehZ5fpHJarM1/3RpibgjBH
dTNPgWXal66aIOExv5MEsEYR0obviWkBZhbb+02LgyQFW/n9m3Xg2WP8Grfyt9NIZhojJ7tZ+pPX
BKBKq/Bug8CT6H1QVUad+t0oBT4w1PeOnYfElSFSYI9uszhRK8G0QNkDKih65zOcDKO1sdc7ZOi5
4nAKWO8GcDvkh94a+O/S6rK35CeVp5f2jz4cVlAxtgYlidvLDDSWOF6qv/0YTq0Pk0adch+EJrBv
arSernC7EUVEqxu3xbH54/LcualuWk9QJhpqJlmNE7QV+M90vO4UBPcKw7jXgDLoi+O4OGeh9Y1t
20bEZe4UvQJfWf6uQF+chrcQFjI1Qu8Q7J94qKSQN8d+SaEnmwxf9DN+OndijlCuPu3cjOVsGOsF
fYnI6HhKXtdxYMn5Xg==
`protect end_protected
