-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZaRAfaRrDRZWwbSSJR3MO0uMIgAsc3VVnVSpvuZ9N5oWJuPAOhDwmsRbzPaoGcORXRC38dYu2oeI
Y2Cku6blTkEvJqpgbpqArWP+TwMujSd3so/nJgTy4OCk/t8m+JNGZtFtde3F+p1qDoIcqtBwIWWn
eWueCn8H8Drw+mHK4l1QWpbHxdegU32+XQMmwsEd/vAwvdg5KZZOzNOalNV2FW2fl9uuyERDIGgS
xiTA8G6msBIswmSyaVm3GfbAgOP6Nl05JFBifudnyfIkH4Pe4mtFDYMavD8uYTbfgJ2IXZvnKBuK
RN810xUws+/WCM6NyH79wrV8DzDCcyGoBmQENA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
51SJWERphwVb1H79npU86s923du3K9anPFbF+7/A7wzqPPcnaHv8pc9BSvzZLJqoUhPv57g+77AJ
roGw4JE66b6cVFzEimJM2xAoKsmmmIUMbs1XzuGdvKj4UVlPp55i2uOQj44kCqy1zWpZtucVXOZZ
eExubmSsWYEx6Nblzt7Aq3KZ0yFYjnsAKw/wayLgQ0gzTw3YWpJm+RRlsJauaNbl7nFfRkkbfLFC
1GdUAHpDvupU13cq1kVvPTZzo9rVkphpARY1Em6dp9Su+DnZvLOBp/ZTSO9ecKV/8Lt3p3O+bNXI
HF6yTsAYCDvSPEG3iTdSj8YIlTlHEpfplRLVFqS5ThzSfrbYwzb8L8sJ7XVXSfW/TJZm0K93C8XI
Sks+V25ZMwzL2+GzpZKVNoOViNfvywvIDmU9Ue6bvyfvWPzx0sLwyqalDX6JujpY97UMDcBkgoFc
IzkxMDC/JeEm7BLK9eLFa1neCyIovtFVsJrMxDAAyyrGQGStuza7amvjEDR6ADCk8vXWRVOKIaUw
zRlNld8njf86sKviffgyKC+nNuA19FqRZ1TLR6ml0AQRyebswud3TtW9v/db8ACe9S+DkNtCIrie
/mo7spioYIiT3lhsASLszwvCBI6C1INg4nWIcpTjAYD7ju0HfqT7DZvebhgsQgxeY9PE2xqXwfl8
mD25pqtt/ben+C3SwCDN3K6p7OzAEgTtHoiwJXPPJ1oIB4z/L9T16wGX109KC0IHGLI6i3wkjxEC
VtOYXzgSgSU4N3k+YnqQTD86jj9bXaJfxYJ0ADfBEwosiJgGxOsLg4gXRLLiyTnlj49o05nfsaaZ
8S6zNd/LDWEkP+6iCPI1GThk0m0/uVWOpWQVPOegTw3vkxckNy23x86nJWlHGVIUt5pmUNuo7i7Y
Z2sCG904oF1OadZkAxcKv+/7fI3AhYm5EB2fkRlnB8s++F1PrmTgQiLIQrdgPxzMM+t1sW1Dz+LK
QmJqz0MDB6vetg5d6IafexgNnQxTxINosmGbVpH8wt+CFDk4xjwMJ7WQQ+0ZqGaGkZfjpcqUcP5Q
hPCGWIkCQBUB2xbMrCAWDKSy7rp7vJnDwN6o91L5xknLItaDQWh/b3aSsD4/AG3PB6aKZnW5z0qG
QMU7Kx/vR3l0lZG9Inmaa1halO0PEjUB7DpJu1zdazkTzuqOYgNvBG7KrZNKiVmfXyU5zJsceXdn
9/2jvSvQW5WOyOryQMLebNJw3xl8EbypMsvK10N4hN54bZxiubzK7gOWBFNC4omk8VdORjfhn8cs
WVJqrGs8vVKwFhfPVOhL7DsDu+OBL0l0XjrFZwc70q4rHJwoObDdEmTI+zS/Zg2iYzfgNXE8W+JG
eOl8U7IwDbc6OTk557jEkuFWxIfN7LWahsnngCihTegWcBDWcDJyjR1mJw6c7pROINm8EPexR+EQ
1361+WjqgllchOkPxcDVq+Dtr1O6JLcGEP08LfL41/0WErjV4WWtlFh0uYT22MLF7D/9jH3uZbEM
XhvRIVBvd1SULxl0PDGbU5EcQpzqwe9FwCtfPyxJ/j2V6cOsb2xE7uf41N0DaQuSk8EVxMUYNUrx
G2UUG4IGvHPh/D/Wg6tpDdtTFX0TgEArFpeNHye2vcxzN3C1fkEre4pk2TYvntDlcPDnG87HRR2O
QgCjyZ/rmUQBCWUt63kAhPac7cBLmcrRp9oB485fMRasiXFYDEZhWwC0pX5FwPun4MKOfan6MiWc
4H+kZTFdpFAON69d71AiwcdthaWgGoLYDc6ZYHkWyJEfPf3GvuH56OLbgtEL17Of85Gh+suRFYw+
n0p2I3IPlOErrpwkD8+Wepu9Pp1P3HZyZi1FG+MwnfaIx1djUcxuxMWYTmF+ic5TfQtatW+/yO5M
1pm9FKBAfiE3aoOKZu3LOzNunaQ5QUtbPN34cpKUViNnCj84fRVkcnaNpJiCWXwW++HKwF+xSCY4
qOpZdeACp1ThAfXqwFfQeuqconSq4VCDFHEIydCvrHG2pfhQLXDgsFq8BWhGS84zbqD63LKpNPEe
BVcYJ03VdlWBttFDtuZi5Rl1E25YlFqQ1rd6b8v+dwV5tUVSKiZfvUyMyzWyVMC4nT+jWnRWTEa2
p4oURhpBqKgqugySRyh9GOSOR8vqtxj1p8z/OhojLs25gRekooc9zweHbrgVTXU2p5S9p2kca9ym
6FUj2/YcgBrgM+hKy0WZ3lZD9tFp+S7q2laoyFHb9GnRXPFNoMQQH/eqPFwY3Vtw+Hqg8F59Ysix
LHXftZ8qZ5i22AG6366WDChMQYN62iuJX2GPNlKLBhWMhCmZP4udtvUBGEG9TRTC/uwaXOCaYHRM
ZzyoZEg0X2QVYoLk2ggM0rJS3Cv+uVgb4lejUw8mQEFyRnSLNDl63rk9C31IXvpWh9vE7YHP+wPk
L7POMf1Ar2GTYPtZRbxmjz0xk3355scTRw/zryLemtsfjF6uwbnIXjRWD0hnKqoe6CpUlOIJkgED
BHl2q3B+vAo3jpIRPG8Fv0mq7q+mlFLBLZdMtsDIrnt5S99IGDxEdxAO/WLSD86tCDWT0gz9ZzzA
YOGwhhY3btc7L/uWiAm/Hc25By7rsP0c390RADkKAMCE12fu6w+RAra2zcpCiRsDwAnpSIYRenU7
PCpGIQSBAX+ReAmR14Z2tzQjygNWIYfHpXd33KZgwJO+hoah/B8kSziknYU4RPCDlbm7rHEAbvRu
JN8TOTykyKB/sNwt1keNHC9Zq37KisCwf8g7i5rcj5jUZ8Ouwgfz1QkEJXRyPfzaeYZ3GikMd1N1
U8t7IFlW0ZPVdQe3E4aGKf3c1bP8HhmTnhjfXwDxBZDrgZ80Vl3O+J426YnZXQOgJg272f5bGmIC
qXAy561uBYmo9ySVUE0GPvhcNDrEpZcVLJf7LmUhXONJ/vSnzmTl9VDJWPpGFTHxG8EEP1QB3Vca
1jAbGWWuj3Vznw9JMoNEsfxb3/NA1sTv5og5Bjg8JO3KNXCW2B15DqrVX/X47PIRMKhfbper3Nx5
Mz0/EfpoB/R9BL+BqvHrR5a9C5kYaipmApzqGaBV/5zSNY4WuYjjHsZ/Q+mza0tUv1vzFw3po8K3
0+fnBTjUGb8DsIiXzd69r1YfMBV4pxQHU/3pLQSY1VCMNLdYiuDbAJ7uTCH6K6nAXXnysRtFcPGO
6EmeFsY9j7ym2tE41o6pLIun/iTTE5M2ye9KVGO1bqlOxptW/GDYy+ACby7j/iCVzpSwHs1LOzeb
wRPeD//Xh0Tyu/+OXF624OK9m/WALhgODiJejPFhFKeZidksYybDFGo8BfmNqjbMHhWlE0yEjntz
/EMt/Ct9wLbTLnqVECR9h6dCuk/fxZIji++Mod6l8oEDrg/yMhjGtG8a1gcGW1arEII+smMLFMia
oJep1b/nz/yQkRRQSA2V2isebIrUzQJK7jcRaC4qQ6TrBTSsLsooV9WtggqfE45nk0YjLAOg+5Ga
IICYLvLYxSTUtECQ/WAEt7hOSFqKvagdnx359/56Zi142KqsPR/SV7IEt4UAPiip8cpDjpKsk8Yj
3t0XzASBET3P6l7ElhYAjiOeck/8/Vv8VOcg52TfSbCju6NLNG1MHnEFEigqQZ+FQiRXZspW9fqF
wmt0QGBa3dSkRVOkeLwGSwGTPwUF5Z80By9MrSTva4DRgO8A8ow1DBGw0ZZQyw24iLVFDRCgTw+u
tbbu+oEYqswkbR6kHkS07Q9Cvh/uX8fazJzsQc49+vbTgu+0Ine2pFzmj/EicJr0LxtTNH+vE6aZ
ymk6AjPxNmfBHSHetlG70ftvu1tMjROeeDobmk+/+dYGtz6gZTFYOJkpbDw1AevCEmBFbp+TI7vh
nb9UpPwSBp1Cy3MGoRMtnwnBEKNPHQe/ON7//COsdO0XT69ukPspyvcLI5TSFhBmW3pvWWHfP0ua
WNZqK6xXtaQHDVjMdW2lge71NoZnC958beoKq6Nkx+KtdlgHHe7JnO1Xf8LyKONorUIz+4QT6ATz
iL8799dgfhDininkLzy9xkYw0Jpz22fjgGOCpU7xrtS+NDt1HG1eZQKr4PkNLDGNvU8Ch76DEVrY
d5VrtDR1lE9gMCwvOeN9qnbVzazom+kdYopDZPJGDaYTakDbOqzIZaODM2AawltTBqr738M69Ron
MkZA4dBYDve9mDMICpdcr5tUwRMW9Ij3V76OpkeusvvB1xJ29eYK774RVNa8caEu25Guu3kLUC3u
NJq433tRxTjGC+EKpK8+jPXSXwKhtfQ+U6LvBysdVy6J5nEs0sU7VnMKzbiAvxS+kTfZYDADJnH5
9zICeH8lzGlpCkmEcnqI6+2KqO1y8tcFk5ftqA8byMgWVJvHKdLnSvVpYYTihVJ9YzHCsyS9JnmX
/DJlQs7fPcQ6ECqkP3GttYEYpLvDTwNWqyDshchtdkxqVPLthiUXzoDNhCE64lwzZnXu9IS6IY2E
GNPxntATG5cuq7Y+DtUxtFOr8MmnmxzhZndEnG+WUOgixYunXAOyxY5znFdgVyTvfIa4nJzLwwJe
loAK7LziN+1hRTSnbIV0awxUvtJNUzAPzd1c3d0VjpvMhfDbrDcLkVhDnpPvBLJH8vWS68ZWZmKU
rm40+Us47NCfBivRGZsiBN7/7u2Z7nx/8BE9g0gEEqz0wPOh2lmw37KwtgLaip/8td22XSmdW2MW
q5XxEBu7LmHLh3QXsxUVBXac9+JJQtxvN+sZITnXqajnX22rjWOG0OZPZDAn9yoCpGBpA4kBnHK7
IlCVYEBHyr0X0mUDv4TAht68H2d2Aa5T/aKdL3e2qYxpcnb0Dx/nF3Oyy/AtsdNU98MltHSWs4Io
Fp+3LBXsZjgvvbornggWuN3MUqHKB1rAHOg3YNTM+q0IF0TAhxLkH9zdDp06V1jIyrtcuB78kKbi
a1i1Py27zCUwWr1ig4KdW0OPdG/doaRvicV26UGRE4aWlco8lwg4lv1xcA+XZN55HnYIfGUmbkQX
c9Fu5jZPjPjhQLfKkX0xCst2W3P19NIJzT2tSKa+YV/3PdWqhUuYyFfEt0UM6s/aklW6iHvo3g1q
uVSnJg1psQwa7wbS81ktp3XTjCaULlK6LkYP2undCA6XndALXtD+ctxLFCl9HR/Y1UbnQQ65pzBD
SPg+7IHFUg7oUXVh2DLxgmPehqHOc1IQalm1T2/yQsqioKP2wpIwNaNNBesOuaz86clonJXIW1jv
lp2D8f6ql+iSwoFBbn/+q4+YCMCTuIJOeBLdb9A29oH5KMLyJZJYBRuuuTLlHzcwPrGvJipkI9uy
VKJ4CL6hg7zeF96xR01/1LF5uTf1VSD8sA4Moksc3xVFA7G70sHihLgpPOx9XfMxrgsBr//odK4D
EsImpNhjwZzN2YQCvfqixdaDcTBeIlaUxav6WdRbfLaz3tcFvBMJF203cSIFPfOrtQqixW/ARBYT
uznetNgoSNoxECauSMgJ1uwczkkDsEOSPMGTui6Wg8j+sGg5FB4/h1niWq/tABv0ncQbQTRXafV3
8Xb+c4X/h7/DpqnMXTL8bjos+wgt5m0LhHt+l/71C7xh86khGHhVSyaH0Ic72lsrzKSig/sZLy9H
Xkf1e1QnMQY6s+0AVxSW/V26AIL5aB0/N6akQIX9llW679+hJOlNobEYBLoivPFlmQoixgUqMtZG
sxlkM1VjHo8A7QxHNAQIAVaijJioziSgeu1Lu66GIxWPRNEKReVCQI4ZkyYgdkx6cKvXM+khH48B
qpi5pgmyYi6PPnS/mpL+z73tW46W1NBEQe9AEbkUy/WyFHMJ1p+DSyHT4rEwDN6ru8uP8Nc/7gtG
pP/nFlDawCEL5aUJkvMl7XtHWSGTaQoVQa5eeZ6nosKHNlBJb76sAgICyWvx/Uml9wtxCU4oLcKc
w60ZYLD2UOh9NVB5oqw+LJGCv8045khtYxFBhQDmCGrBcu0YlZMtoylelIvjbs6EP7ZBpsEZ/I/F
plpy6237zN6PBGubUt3yYKjDqnOgl4UdCFYGVrYDL7ec3kjE2jToEy7RH7E8RSog8cdYttopkgpP
yFKMwEtJ4k3T63QzjGFLhzXzZro+H/SU8OAYuiyd+QDCwm9KHMS3dUP2aacOE/ulgwSo4cytypcM
VAMTOUh/bqvK/SbHFOoXpKCwnL19SdN9aMdbbGL4N22RubHvimwV+gYkHIxBlCpud2hT2znxhVP3
COj6pbXA6JcxFlBSQ0NrnUBMnHBxOPLEq8VJadWJkRbydoXQahR91gotJ1WmonyLoQkhaD/QCfhQ
LgIvfLZfG09LlMlQuGqZYB8d3x9RsUMN86v5v4PJTZNLOrUACO79DwytrNrukWWE0zXkg+qCk257
3J8O5jVdfVSs2thJLAOU6dhZiHGqSdatGm0ZTcbtpefRP0zPs2RyP84FvoNmBdytfkLwm0YS70vb
NdzcZI8HXyw3vvfUECeLT8aZoxKlrVaiissjPl20cFygNfnqPs1dEeUnq+TEJotl1GVtJsR+5Oti
H5/czqPE5uuNRQ2CD0A/7gnchfBFca2qJoI0Gp0a8IeJfhP4QzKwtJvPHOo+zHLD5rf19qbBeXWF
0tUodfnMwH4c8VpXoRSVNXzJF+jMRByANdpdJ8r6X/Z3xD2wb0biiJIO008qtObts9iWySHKi7oa
RQ2YBjfR/kwtkagwpaRCVp11ZLHtceNyNHvwAYHHdTf76nj1Kmdbb6JOyUJI3536TsDyYfGeSriX
e6sWqRlN92AjRzCXZT3kQV9UsygyuiPLC2mW6Vu0CeQKGsQe/k8/NPCVQ4XaA6M19nxmoCD0sGav
7wJYevEYIFd5+MroBFulPSDYR/7W51viVSoHzgZmzyzrRwiA21sHld7oS4qiNE5EsFXml1xXZXxU
sFW6ygZsC9ZJViQ5DsFrviu9UOdczre2bbFG/ikIRQ+xZOr2HPbr2RIgM+1sNPrkz7bXEDVQLP12
s5+h93uT5O+BdYguflGnNJk0eDuYey2UDa8VOQLcactezBFaa6MktYccOmNsyw2YFAzO4p/L/Sbk
hA5cTTA2oXlMg/29aJeiJeCSCs/U7Wyi2RskBLB00zUYeTyQDn2fAI2sO/aCjyDE+YnxXTUNadir
OdL/Rv8F/snpTELQFKGkQxZibHdtvpTVckpeDYYoHaT46Ky2BPzEgMPTE4/ClgELvvQzCwPKR2T4
AQw9NraD9Z3GSfRTowBYs/vYVsnixDxPgT/4mAwJQwbhuf6wfbteeoqvtFRuOJe054w/NiHk8f1/
/QTPDPGo4duftgTcWPXDbtIH6/+mZ7H4XSfROUwBxOG6Be/MiOijbBgdox6/8O0mpHacgAh7q+Ka
kdcoQXTJMOA7lfXBmbRD8wiLS9dlfeQLyETeyvDcVHN8QwKJFKvxcGhlJ1sSfA7amoy5xhVW/08Y
bg/QbEUEZ1miwuIfJP0XctLBZW+rEu/UdYBTPbTUotx6gyK7TEtna6dMah3XDB265MhKl+t8ahCx
by3Aom5YLv1d7lTeBCTlm6T5FlGzBahuznFRDgj0/9UugsQsKvmxJGhDqAzLY+DA4eu0JuOcxfxx
AcEg1AdIGFz4qDfJTXXK3rGjFvekrpkfmIJemvBybyCqoTgUjXcT4lrfxjRUKJY1jCbdSPTHxKpT
HqhzOua9rM+YubQyPWvf1I/QEePqfPRDZpmh2FQI/mWO8DpT0L0NGW2rsB7IHuREK/57lAGBXKKO
Pw7T+oDqS1hxk+Svk79Zq1V3cOpp9pMCSxTPaWiJQDCr4KnNIC42dZNak31vzFoIw5MHcox+XVy+
KMRXJ6ClKFpdQ13bjCeQxN6DSGZ5gCqldequTcyUl5d8zSH3EBLTl9qvL7G08jblsKqI1fwxjf45
XuByht9O1NzufVLjQMq6Ik8GG1vX3rxOR9DAnnW9Ztf0DqQ1RFdvjqfJ27wIdQ86r1To6MP/iqAf
2u3++KQsNlDW8/A/uL1Sp9rFfjPMNHVyFavKX8LrRTxLLiEpFaIsh3SiFRKSpDhYtL00aA9wyHdB
DdxO8GvciLZIeCHkGKsZVCh9AzqBQ+t3z1iTsHhBMORs5/tgCIOFtxqM7zIXXBB4iU61pGq1zx4e
cdAb5ugeE/GwWXvTjz8DPveEnq0xSr4nni0+tJaifDtw1mFCScuf9RKuAORXxBw5oJXhdMiW0VVx
Nfnxi9+jc20SV3apttLEsbTfiOUZFN32p1+q7CMjlsriMOve8Wj4tmmkJNGlYfMuagd+d98uVm/z
03qbO0JprpQDJwrOydKfJXIcfdCatmEyDgyEUnpJWT0LX6EEs4283FjE4yXZYr/FTQEnC+HT02GA
H1hXntw6cbERTeYe/7/HeFi6pL2LOm5re/NWUUUT2CQiVkTSWoxYPxm44Ua9rzFd5NijPw4UxiJh
G/Qh9C44D/GmLHLK0fw9wAjzVY2846+0086mvgQ970AfGg6/dAS/6msOSVs9br+muo38ncwIrxB5
wq1lLoluZUEJadrvOKl6Md/s0HIo/tZJYO4fkzt9rV/4sjHxVEVq7jsuW0ZyO8K6fwna0XuudDFh
rhCyWaaXolBVago/LVHg2aHik91Lw7QeDgkyhwNLpVY2OtLWJk2wfRIFuQqjDmP3mlA4qkl4Kh9p
gK2hP9OSGcBBNBnHNmCHmloHuw7VYzb/3dGbmZEBnSl0J0v/g/FcnR79WJTeIsaD7WuSxcFrUkCU
W6AKEkzNswhiUaV7ecfpT6kkEQTl/09j3ihe4jR+TsVcx54dUDU3PmiRNiqqsOwK+N+q98Nj+6CS
mM8ctbyd5knny93pHve9BXwG8i+LYLku+l/mI7J3nNjL9W/5EWB2zsEK767H3e/YOPCRotL7artl
HVGjVWNwZq31mL1pvbne6A+ntY35E8sTPW252JbiKWdNPdxDUKwHkfKpZh0dh1ZvbbX4NNwZBF5Q
a63PI22MT0CyDgbhlzN4yXvSGAaFDPG4fhbUF5fDS6ejqV+6+aZKdqh5NFUwAMWzcwTBcsM4tyqx
WLlDDWUEOYNNmoIuh0NMil+ZY0itc5gJwaMjJ2QWx0xK8/NlGB4/mrAj/ZbzxbD87aTpsBwZVkg/
6ZjS5bOl+0BFYNGDbsenRszXtgtwKRgKGGm1CPKs9O9NokbkjvaqcoFdTYEIjrpEY73XReXtqngC
ShuIORtg/XjZgapD74Ebhs5a0Bv9/eJRdvmxE8cc9Hau+FRKY03qWSr3C9o9C2dIYPbQkAQpxQlB
zrzE2cGL2jWUesEGLmLpH89K8doEEQBUaZGqthQA5zYMerZaBFPyaoz3HnHsJsQxyXHyaojd9XFK
GUyzYrlZ+TONzakBgVHpuuzfs9bGelZ0KiHDKPqICzVgmWCQ5TiXlh+dXxIRDG2jRR7v3uhOShUJ
/jsfjg8IjqKZJR/brUrIYlCs4UDPpNy+jbwu8LLmHVWd0JUQ/cjcvJ924euE02iYdWtYm1UV556F
3kQW5A9H4TmbraEsaU4QJc7tLmH5KlUIrVayuBWS1HPwNPwa9OKTKMdiqmeDv/WXbEwcrdKB2Owh
mLp6t+I25ojRJ9L+r6KvtLuYRZnJwwcPNWHWAiB/Vf3Nt8sTpvi+2PTkSBFTroB9GFqEG6QFk085
3CflGfCfGkTJ6RnQkRjuE+2HDZ9xq8jDXpvEjm7cQw4xH7AtnDuZUMmujACwD4KmY94ESQlJX1Vk
NkkjwyFYjw3iH77Zgk5YwgniyX4GSZP6d+peWfiBJ/BjmK0oXLJot8b/PPqyV0IKyLB/4jFrnC5m
uV0juMu90MjlugpE4Fyibbs4Tv6wYhQkxMseSpqTAC2PnTJRMHIHXRM1XA3wpZqdUK1Qh5Q4bcuD
ZmbDkLKjYW0f5AJJRH/ayY7kTdWvtg9fCf3G8pYXJPR49Ze6J7PxJs0MYe3fUmzSyJfaMDRfhvZu
YBi+RmNs1lX9Xnud3RxUf1dTikbYbS/T593NSvk6m/GF0M4Yd216kSwCkxZRGOffzG+h2X96VrRr
8JuD9+Uk6XGrGyWvsrwMG+tBAm+z6fYr9nggb68vhweBL4kSdlwc9T3JgxKbYVlhZ0EwwgWf/8xj
eMqu8uVYx+x5zIvEHv8OgJbNpFNnRNIQj+TGIlhATphyD9s3lgn35ZNe01ATcjzIjtZ1QEVZFn0T
xO/ANOWfxJdv2aKd51XkvgBm6cZMPffUN69NiSWVmoYf6Fltqk5DTPuFHCcK/EdDUtFbtPnfqlTp
TAWCk+LejPqj9aEURowADZ4+ft807oNCXrHRiFqTQJVP624tO7tihlmz5GFc/WjcA1D1m2ZkWo7X
ArtHTJIjeiHNmgA9jyppSPKGn4Cu3qbRNXsUhFxa/Lul2o/mb9ZwSpn5bmjP3+VD+sCDTw4A50J2
hK9OL7Qxosr6xQ8IQRXJ0F76eiIqZSnF67cZTaPRsrz9GO+DSGqAVBV/MOetSuRsTQalU01WAgIq
jTHI0f0zn5U/HcDduzy3mtlQ0taZeNs+huyIlHIkGTu+TylpFWO0x7yHIAabDFh/ZwTEjpSX6mPf
rBgJmSpE2xwoSWNuqqBwN+/Y3G0/RDSegMXdkNz9p2uJwf2E0U4WAbWlyH1FigVV7q3je2U1NX95
c+ar1ke3XFZ7EXihCQpUYVEelRqCMGc7TOLYBvOjHNrEppKEbq4cXB2Cq112kx5A+ohrVlBxhgw4
biFHof59H+yQf2Utdtzj4lvxoWcGZlC9bFefG/75ptY6LjzEwLVHhK0UyPwQ8JWiQixe5TQxQEjU
MyCcLwhlrE51OZkmtK0XxZiPTFW8kK0V22xjuExox7bc5lUQuHUa2Mh1l3e8BEnezbggalM0b+ec
ccptnFz2izebPJkxPD86xtjPlhtqcJZH7Bsj5HTfiY8JxFuEpGtzFhT1MAX88dYFm0rwzHLP6bZt
KV8xRr0qtBuPHaPqnj77wN4WyBzsRg1dJAD21sqx+b6dMOxW0O7bmG7slUhKYXct9VbHIuexWI3L
5GVdj4jOXrJ3Wxgl9M00wzJ7OOJDNCnS/iNOz5QrFuCpQWoeEbf1iBSMwslZj2avWoOiQNl/A3ZE
rMxK/m+e0hJ+laL3Piohx3HnEzWfJ/gb/80gPicR/WtlxI3ErCzN6aME9ck8Itkd6L4nsZs4suPj
YfE2VHGqsZ2pSe9x8EcH+8MASEj71ikw35kVlrGSyn5PJf1bwYPuhx/V2u3YtYS7PynqBAxhHA1X
zxZ7X1D8zLVtwGzEKBZDCPCbnV5nwNjAxTkcRSB2Dfz1kH1YMGMdZltSVYlA3Z33tD2STmmz5dfK
EqJTezUy9r+p7m0QcvTCuMA7LVyfnSpIFHHwguqPwrxKf5gOucu0MinIX/97fSjmXzti2saR9bLz
rgmfNk+jIkUODx2Uatb9XBLMN2Tz3vQlIVeHlDibz6sv3zb3D0K2AzNNbEIPxUX2vKn5KgleCSAk
UlcM803juJobUsfK8EzrUWpRI8oVhVDcyrEgdKql683WU3O0f73N2Al4oRrrRNdCnKY3ZR1k+W7X
rejzC7MnIsaGvaI2V2zMxGRn7dT2wp8CbN6mNHNMeyMWH3gJ5pFZPvcomsRBM9bGICgr8RXncJBo
Fxf6sOYp1AIk5+E82VkphNRB6LidOR193Z0eXlHRWZmHuKNB/BaeDqYRHZwmHZZZLhSpgmBNbicY
K+77yMxd2I188bjlLwFhXPi4Xtj/2n3dEfB7bACclWQLdV2O0IwS/UTx8WNWbrafMVF1TEm3aN8s
URBlUv7MK24V276idMkgTZEUt5Jfu4/JlT/CtVt51flHQasOIbvZVqv0eJj0PyJj2A+zfv7BcQYr
FSv/Ieeq264fMCuUrNkyHbtPFBPXlLOl+b1B0SBe9PLiIypJUigbyvLHes/t51nnFDLJjaXWXuwm
V7cOjvwdtebcHNAPEnL4Z9W7HoFvEfYBaIgObMtkwoTLhL7nElemP8+LMrpUxRB9f0cs/Wo25kn0
whVJgMv4zP/Ihg5aqdHNz9wO9ZWiB3VhKntXDo2quSFEM/MsXT3IUZlt+8mKQAb40Nq/TPEmE5Y2
0nm5lhzmI+2A43mA1f8iXIzvT1BmexKNiJ/Xs1dVh18h1Yrp6ev4Uz2PTYLq++htCLh3Z4csLVOh
p6qqvS/VAsrMBrAcP6Tl6BCi7M6PEvBdJMsdMpQZmHe3TlBiteDnMsnQ6NyNtFXNX5o01+976Pt7
A1iI6xLo/OY37NNuMqKPDv696FUlh1Qa6gftELt2aE0ti0J/UpiUGdJ5JkFSLlv0myAPoUEOgMLg
OlAqQPrckhDI8vyRe75p9RJt1nzBomwqi4PL8iyyiPnbf4538Wh5fqFS3NZG8z8KNMomnIzSWpg3
MAJRDGf4ciVEznCELRy+yhG52FdH2f9VHguzMwEaMmxvbRRjb5o8hO4nQQH1k0DFbqtqpZmgl22N
Q4NFldv4omR29w/jdUqwQv0CL+rI/NWvY+Qz0HxnYhZAElL4fryeksg/NiokMT2g4AZFC3hET4Dy
fNzG4NVY1Ji4s+/pxZTL51nh9tWIKl/iXMFhtgD/SIkVPlo7tYoMxjj87UlXcObXwGvbYjITOeme
IIH3fwllxefF9I79SNDGBdpIRavpqG4mrzFFKOLxrbWMe5wYXuS3e9x/sQmUB3N8o08Y0b45x9EZ
EKQbweOJbOJCclzrF1uHFJCNIx/1IAPGa5qLSisEfd9vDCQlsITPL9ARS4ScpjT3an1j0dYZhHD1
kwM5tPMwu5SUgDe+uU7RVOtSKVdU64BEi5ilZ0MhWdq3+yBKqfFUZWoNlARHNb79yFXydi/CfMYa
56Hdx1y1LGguftKhcz+sGjk66wmH+WQtPJfynuk19L58PVy+omyuCkAcEfwMsnMOqaHWfoIcRkVA
vtW5QRNfeJozr+rvz0dTi/n9XpITPPC5fSM3Sw/0JiWr7EwyPMizJxNfiom33JrKfMpEGYVniwKi
KbpmAHa4xgAWqXayVkjdrbW5fB9la8w6Bis56dRaXVW3LkE5OilFHltmUqJZcqguH23QA9dm2cP+
GSKhVJDKUH5ZVU3HwLsMjVy8FqLUKMRZ2hNqysXUH3ZQfOPaOHC6M6R8yUJbCUYjIBVq5pKDYH+c
8u1q8uqlv7FUd0nYHawwbT5ihohLPRZ1MDImjIxOU2SLUL6xgRZbFVOD09ThQelXfL2Li4YtoSSi
tydv0mRjwGGwUTjqQgaqQLWjw/NKMfMmj8AHmcnothgu4TrN4lqx6BHCFxSruN2BNdGrFcmSMl3Q
oh1p3ZageeeHP/9cKviuHZoIeLLSymTVyN7bzdc03JfiG+tx7mnGGj+UsN7e4Crgn6elFVdh1HJO
9fSt/Y8vkeP2FjHBDnJLFsXpKxJBWviqAgAuY0mZ73+FZqFlLDGeSf1teAMUrbtMS3vaYyGn/MIf
xRZ5JsSUtLKXRwjfiNzRIu1VtNS7zlbp4hoic+7ZvNz9tLv6exWZG/6H90wwvlR6HntfvRSshTo8
uID1zM/le9hBMw2LjuD9Dezd2nb3f9xzRaSfdeE0VSvEm2XV7Xi1rVcdBLYw8/GwJRe3PIxAokFI
g0sSkrgo8pGShOP8/KZs2fgVrWJgbV6nj3weNmrwpSJFj7FRL8Sr2eCaCDJ2LYnjAdPYyJNWc248
5Ij6mH6+xHPia7c+LxEVzUNDhsLDcuOhcofdVDYzunlRpM9irMvxTtN3g7jxCTokpVQ+Ie3UcghP
BAIeYj5g+yRUKsmTPyu/fwTsBpDbWmvUxuItGonIqeANzZCmFnh0tyPml3vM6umW+ygSBSRdNCeq
h/dUBvOk2dzyEehZCNHBYVt9Tf22HuJ57AMeimLnVEeuRRFgcXjeyornotSEiTR7ALdgzYBfERkI
7ZKSZjduA8WNWuDipU+0ckLH6sozT3hjZTq9pfJjFNihrWdWlO839s8CbSNPV6mKuv21RXnFVaF/
dNNVaX9MO3y03Ia08praRnNiAi8MNHuQHY2wyIsFaGqlPocwkl8CkStUH8raOQdetukVM6H6rGWl
sbpkl/ONLhMKXZ6uOTFG/np+tyv/tooz8qG0mcEGXL3MbbxU1T+Zv9ai9G64tv4JcnJpx7I9a6KJ
VzRQuzS84qiK4S3cEmNIfik7flfmVo8Y0I23JMqRkaONCza1/dCvXo90wmX0OcsD4Y6gPHIiyx3f
DYOHyfYky/urAl4CqjkMEOHjWibDMGWDiXSoFwPq0Y7SzuMK6fjn70qqwEtB7Gv6oluwaf/TFbtJ
Qb0Kxt5BepKa+TWvrV4mIvbh0PfMO0laj+1XmsulhoRbiPSMeze/Zq28iyin3OfoI35rwrzVpqgY
IsOPg3UGgQQxD70FZJsrbDLZIc/K8LoPPg5ikRvgFQptnkKZ2Bu+b+NpvyRAfndXaZFYznaUPDCs
/H2su8VxyzHQfkDfhBdrMELfaq78LiWwmHLqCMnjRwXk5018rkLJQfBwg3rFKAMLDUI1ACjHqdCS
1zcAzA+SS8LdbshaDUeD4V8/wwfVLZU6oCxi7/BZe4+eRBAQwWS107QwJVN53f0sbUvr0NptqhZJ
xOsZV/OYr0xh5vlp9Urew0BF4akBd8x0gDOtn6nbKclloD8apGF5Gn6hkFjnMZnBbfrZTS6KnYoP
LsuFYIsxnFOw+eY2EFWDa3Hs0Zh1OE0KhcNg0BVGq2KegmRK4At7VSimfHEFB+0enyn5zwGXd41P
wsF4JZO8A5g8NERYUYsiptYeSZuKuep+wcqHgD2CRg1MEwWoI89XZlZ86FwxCPkxacvBWRWtSR54
EdLDpziLOj9AW3QCFn5AxaXgnRwpTpohUoqc2KQy/Htt2HYHK5dsQ3AIBqIay3ZeJFmFatjdIGhr
HTqOlLLrjVN6f5eCJYRktt3Q20JYMS1YUjdyyi6bv4g79T7AR9ruEf5mdetSW4YSgHr+G0aRNK8g
C4EbugpLJvJei8a/RQwYC6rAy2msQuaFDhpEoHyEf+dYtQLXy0r91DWxFy9vbRQNhNyAHSSf4zr7
cdzpDzjwnbFeeu7NME6eDNZ4U8MGuIwkilL5cdRCyqPnOjIS+7QuQVipiTtossN1YmDwDQZgJRf4
fZAaCahNwoZNe5+Yu03psPZPAcfy0orJ+H1xY2h6Ao88HyeNHgWkz6MP8bxMqBe7CoTPiaaJ7eN/
uWx452ckehsfN9HpZwThgCYMI/uA3HB/4sLlY/xq0WK+rc9/AQenqF7NKcbFsB1c16XAe9Q50A50
+3sRjNpIwWGkI4CcdRxqfwieiGQLLOHtsAIrJUoZe3X27aJ2cuICT1w8ZRC4bds2FJJELj2jQNMx
QmIizR4QzKUKaTd7P4XXa28EfjxwnRGS57rOgsYfAE0dT25Rt6vluGShV7Fi3lSJ7+WHE2oobpq5
Ib/C9YQhNfxw/ZM8ShVPdm1CMMGuHBgxLPzMP4okY/E5zbUOi15vGGy2jt3yrdMHIt0UQd/6xwi9
HkbLWacmeIeRkK0qsfIrWWw3QUvM2Ilsj9T34odm78xMppxSor/I4RND6tESmb40+wkIkH8YEXtV
IEx3otNx9yccZftJdrfc48H6b3h9SAsWSy/xvvb/z/b9Nm2Z3OFnj674GROilZdTVZxI2eWkjEe2
geGYB5JrFOMWiTZzawyoj/VfD4X0usFwwNbt8jI8G5Lwhc+Ld/QXePoc5BHPNbFQN7HcqiZNHqd/
NFaPHBoaJ2Q5dS07ZkaQF++KIM2SqBCLMl82uQtnckpfrymKT+ymQAXB009bgnMUAIRgqo5VhE3t
bWCimUUa06hC3OBDslx5SNcfSK/KbQtE9W/PQ/WqhoCF7Zq7MXW8u4HLg1ovfz5hOnxLFhMMGiwB
Y5UOrUse8pIJnRHPnsqMLB3mX/hDJU+xwI5aw76XcIAocnH15hI7nZDCyQyw7MuAAO5EmlRgARsz
9dg2c/6UTxSk7N6NCMT9r1vgdrtUyyBHLw2pjxdQN+1zHMepWWNHiUo0kvw52wA0uA0NZ62jtiDT
Kaq9TBqJC3BJq6edo8yajG1c1APgjTT4mMfnhk4CUDLIF0bojFTgQOa6u5/BNs2wapv1gqZff0TP
YGJgk31xCp3hgVl/VqAl9TUYSeYXbdMFN+sREAhnfdLQDDxjR5YKRHWer5yYeNDpWABPLgYyfDFd
ot4Oakh9JkgJSzKbEw7AQUWpS0aQGVdmggAqZ/3GMHELwlpuitxzEeU8dapRrclFuZGfCVPWbK1X
9Zkz0SjuhTzBb3NA0AJkNwuwMRJjzSrT2YxmfDEcF1/tUeA5rEQzqZBOKswGw0lcc5Lvpt/FfOiZ
9W/UMhGVClEeKmhLZZ1KHlijqXeHRu8Z4zwiKTfDV8EDVzv9JoJ8/71dRPnC9foGCTkSa513H+qv
grztnfFnfIWAXE0Az1eAy0mPT2jDqEBU5lrH6Eu/iFxuohvB7drRLQpAusn5QbrEAT8WEkYLT7vP
IvguN7RYr1g9ufLu+ck1IWJR6YQiH0bePtoZoXORWYA0jD7jkLZ4WYseCohOywXL6bJ8rn3KWpfV
BetwJxkZLruxegLXROvndJc8TYJ855HW/J2BPCLpSjIBLsHWc2/UOkPQjS6M5Hh3LcnL8+rOQHUa
PfY4/YdLYAn5dYM5tdpCsRs5odKSCuxLJ/rcyQLqGpqDBwhaas2wgXwFLcTM/TxjBQdga3Q+QN3J
T1gsHnes2ACzbScjHer8ez0xrWxbgeK0BQIU/pZjwLL5o49zOPsJ9o0UeraUX9HcWkuMmgsdY1Q3
ZkcpPpKtM3eipdElnlrbCNA8T/V6qgRkuGrt3jmcZ2mdf6Nqhl2r67wQAfe0KsvoPOe/9AV6mT36
gL6kYPH80KoiikHo7+OhHwNXmX0dX5szyF6gYfIL0s7QG7IPu9BGI0brY7WrZeFyjVZZZR5aWVhV
vCobrQ4avIoMET+cFxgXLV3p3fYFvQ4P4IKS++GKVZmuwQLQYxNeQVWzQylC874zL5K4THIxaJ/S
MD5bEjE4ETg+Yn4IpPNwva2DNdNRPJoPC9RrNNh6tR6KLzLk3U3p76uw60AQcLHho8bi7irxWY5C
jjUnLy1gDdYivPFG/Mckwio8emef7P4qiMPqqolbL8R9T+Reru24O4w6zfOBm9sA611x0au2oEFT
LKBl7isSMB5Nt7lZ7hTdrfnapzWTfPCwwkw6CTLrGnSA9jyS5rutYrOP/kThBHwKJ7gBMGKkXCrU
xxZo/Iptz7BX14SzGURGSuM/wq+JhlNATZdCnmepnmZdQ06Ha+Npf3hanb4qj/+BHxy+7MSDFmVW
p45qcGvpj07I//5iAWiA1w6fiiGduZedTBU3UilDyNjz0UyAMsFfe52wsREQC1etxeY6cQ1w9Xc2
xM2liHEJx4Kh6mltlCFF4sQwa/mk0iu0wuaZS776Bs7QD7QAcsjX9yBQfJ7ef9i+pNxRtelgJL5x
PiWH7mR3GxdKvmr68JlRp+VDTiSKPcRLobOjjkmPI3rw4LhT3aFWYRLllZdFQU0as99D/JHmI9wW
6HyhIPUO06dFTU90iljxT0Ib6hRTCsEH8Pe8bQ3/kyAjJ788BTT0i6KHObDGyKA7CvWModJOjXzl
RRy54TiSerecVwGreOHs2Q7XzZCL03MnVB3illoPHcGjhzfKx0qGcnUd04Gki7Z/DYUZQQcbqw3l
exkrEmebH0ua4Q5CDgHrNPev22ibZKDSpdzlnQrZxbttwrx0xQbTv65GA8CIWXq/0zgN27s5JcuY
Zmk2i9hYjZesmR9k1tOkoiAaMcIedFkXq3NWsakLfSsBxZvtVQXi3vljJ0V6pqps+pW5CySDk3SW
idU3EvZ8FZbfG/NuqnStJUYaY8Z8uPS+sZzx6zKE/j/xsKDDZfLKBQeI6PD7SpBPeRLaSBAnR1Yk
+6V5vgaJ9Ke5X6oF44SRnpxRY457YlWw0zKrba356sUtJ0ogN1BIbzwdlPSrR+g52m9TDtE6s1N7
4oGxgRiD9Rf/ds+FqbyL/yGDvSeSQXhQGO/MK5L83JpVAkPu3InP3PQEDe/rUronu+hxAB3c31+Q
CjoqBfsUcm6l5ICjdpPfTZGFIo2x8DJe4Qi6rMzwsykFiHcYIY2VYCzp1ivxj1N8yM6d/Me264PJ
GQ6E6NYZP4A6lma8O7+bvvlc57d3f33nXx8mNktdCXAFELIEJZcFuWRK6ZLoArTlRbniRJIH2/mC
ZBckx3wJDkMWRC5zwVnqxP2fh2Ms50cOmu93w6QwkalPvHzQppRkVUbDcR9F4EcnpMiMY8+VXnnP
lLYVeQ2btED8GPmMEM/GybqsquHLd41ar/5+ovgQLfwvRZBaN2V//nOKvwbec0imGCxqFWJ0RmW6
AgtSQE2z+Tq2N72hpdFlX6QaV2e1grzSp0XTJyf15uryiW17KT1/AaIqU1GjGAas11dS264be8od
O9JkQ/c5xUaUCy2epvckWU5W0i5tkFUlVTUnOkG8XWO0IrSELkNWk18NgCm/ZZktB4gKnjtK6YFx
vAdtyvHoFcYRDu6b5L+GZqLijtIK3k1Ysznc4rcmV3ALMeoAQlVJdbLzPVi8QSE9c2aot+T4O2kt
AbIlEsSf5ru1N3r1HsWPWvs1MFN/PdxTyUTS1XLQgSJKL4pXC0T6Cqu/xIA25+/0ya0YlX/rO3g2
misag6qNZ4PoMocOrRWvoGvF+54XreAgypOF4hjksOvwgqj5NFBDZzXWUy+7CgBneX00XnTBB2DR
s8zPyHLcloffKErwVJ/a/jrb7/B1+vYt1ADcdtZdoJoCmndOUC3GM1yfdU+sesKlz2ZxZi+R20FQ
1fKLMidudRrVhVHf3CpLmXRjhmINhsv9jtFmjt0VWGJ/4Q/rILdYA8E/DL+adFSo0Xpxa+lnm6f2
IHac9RMF/cn7siJYg3PvcEvel0x9wxDz2mvtLjwrzSr8DkhEhQ+sBbSB6wfNU1o9TNKBgHZ429ZN
20Fo+p9Mf5HyMdZUbYbXZPQbaCUNvdM6ZEN5PDmlQfuxi4QIxqJj08LtEl4UqkD/9IrtclClXq2r
ButNiKYaOJlN4Uedks3NRhPzGKjq2D5Pa5Og3VhLHwpVx8WPDnD/8plfOHJrPOsIUgrgnLaK0g6v
bzKIVc8/TCZwtdzGVKf0OIhxP2j9E9vyZtSHAsaQBwzM8XA+AfCQS7UQIhDRDH88SX+0XUxuvufd
wu+cHb0M8O0sGSCwdrMYthYLc7h0OboMO4Lvp+pbIaMW8fmv+6lv6XH0V4zic/olKCHMBD+yryKF
E5Tgq9JmkXhwXX+TqfdAv4wqUAtJc36FBZPCrEhfKsH1XXT1Tl+D3gNHEveML7UHLO4nSOUc13Mm
EIJiK+ZJb6XMH2v9qCuC4BdSR1NGuPVlWR+TpJBzi3vWw0qp1HRiv0wAWmrgkHq1JzhlYpoSF/Fu
QnNIejkAnG0+XLbCHScayHl7pKWdQOZHPvKbr/VZa5vyMbrHEgxX0Zc/r6o0uiVU/3T0QgDpqkYt
DtI8wXM8CZBzRDTXP2A7aUhvcl/hDSV5+AhTQq3tg0Lx25t5+huUeLDqk37FRI+OMr9VivHYoZaI
VdLS5ZW+akHOINUS4SUoBUhR64fkdeRm/iAfcBxW5NWTL2gdAkEjWXzwxvTTcouQPzeRgPlWpfCx
YbCLiO53w2Kn3ag71TMcHDnn8NQkQEKSgZMw/5OuzkDOK82BLJltpBUjWK+2fqeH8gO/WRZW/pcn
QkFBAt83Mbk6E9iSTuypVBa/1c8kHPt7+M/HChHo5H0DdbX5mhTfevZfIVNtY7ahSshuqACZ+gYG
QpwL1v64bhPsqmEqtFhv0uI0VrVrFxG9VLZF89WTyqkZVWoSZeoZC21K8BPgxOkCi2DRyx9DejdD
lUYqT1K3tZADHdkkxOQoRNoWC9GhPwxoPiJqNmlpZJvYr77bKhc4xk0wuDWdG8/R9/cRXDilheUi
MByLumwtFvJpf2dniD7ipAdGE5z3kRcXky7afBmGdbdIgLZksTr75Ri5e0lVmWsGxQBXrsQQu4NP
7nCiyukSvN9124GAutHPphr/G256OvDC16rgYr6riRXV6dwDFJz9sREbazQt0YiO5g5kJuLrnB3u
KtyO7zgcltK0PCdfgbx8ZLn7FN/09lXo0uefaMakxSofo/oElS6Tu4c/xOWBDEUAPmuzM3mhwELo
N8L2di8dCL3TB8+PgI81KTaOqWIhXoCAkGHl/PEovVKtwsPFoqY1zTC9cs+G1txLrlSkfytQ8TRf
6PCjGs2iDc+SR7Y5THc2UwGSYfwSlGAZqXPoNjZ/T9NIY8+P5xk4Zqth7VlIPIIayNmOYmNyDvjw
HEkCewiiEJYwhOPL49/z/t7PWul8dJFLwKyiexONP2NjMsl+QeKxQLmmdglOpKuGZpf2PsJUuUmA
Eg6dcUa+Zma1CHP7eTto4VlqL97kJp9kILhQEBVEVx2/f6Tf90NTagQofUuVatOuCrxgK3Urgb/y
6/HtCDUJc1+DA39go7ytWMFHgOowvtxgYwiHIU7spDcEpMxqGXZxh9iN+Ig9A1rqeOVz7FqM5DKG
EGlGJM8y4q5o5Y26WTZ1rUnr4sv7HH8o4xvyvHRLqZKtoEFkpfbTzMaZWrvrTxjYfBGkoxg/93y8
0psuvj/3XXjIdtYe9pHxTxyKbd8/2a3vtdZGyuRoLnYgyJmQ6hQq08Yt9q2oHGSRpH++M0HTxX6G
+oXb7WAAcOl75fup/1lBPqg6XUs3DwZkY/bkhzLJooVQ+hfgqwvkeLvHHSjOKkpqsQm5Qw7Pbhyl
GPOToxbvuczqM2bn3So6v7l5DcF8/iAwC6M8FiS6B58YbkSZIBixNYBuhCymJYN2QjQX9MdLO/p5
FMYY7DhCUEaxJRpRoSZPKtROo5a4lGwcRNgYIzv5Ub4CicWdBSTX3Oj9yEEClSjZnqVxgfX3T1Sp
x82BXDwEuZZzC1LPZJdFqnDKWO7IUqErzVlD1ZpdyOScDgY/xIW4RxtEeFjwzG7iIpn8kpYfu1sl
1XBDrgHYjms/5jSDFHea00hBds0f2MRDa5IrWDe7JhZF3Hooamz8aHnsNw9RgqMcnENnc/2Unpj3
584jAmJbcNcMxvHUTpXsPOd+Lme3iN/JWG+76jlugAQD+01sQfLFKWrPU0uUd6vaPHO2OPtQAMDd
Opf7sZ7iz6eHdj8TcrvVz7mGbu693rtxzkxvv99P2VgisPrXNa4LZ0sJVpMccCgA4QMOmiT+wbp3
lF/OQBxFcdy4idyXJf3KaU6FX7Hu2oPAOgb0fmhQSIYJ+tXm/rqDYsQKMozuQ5BhhrNsmp4UihV+
Fzciscf556DJqfqE/z1Td459dC3vaTaaIDas8AkV6ilSUG58KEDLNjcZZAj7budpQ6nYhzNUdwne
krwHfe3wMRReWkJ8psf32j5R3AkBkVkxJutgHOJZM7n4tWqjFfAVx0FDUbEV0rGc1CRcPvupbj3t
JvlhrQIXhSKhkUGMcbo10dHdq355Z5dsKIOobP/e0DTRkksxCEs2Zl9idx59Zj4GMUNsUWBQsjHo
A7gmlnMAeE2Ag0Hk3OJgi1K3uddj7uqUN+39l/VzOHHh/ASstVJ+cOYxKdEwSzahdc4uJsH2YfCQ
DHcGSSu8LINC9XzgKoT9onOY5797I5C1405zjiKurzj3jrzYWs0C132MFcgxlLiz9sPpKSUeLD5u
YwYJxEn8nQ/natv9BqTAlDj9XweE/fK6pFC46ALzxfKe07oKlLwShQ+PlPwCpjNPBTOxYjViB8Tg
MckIhsr4flYfYcCnl9a5/KH+FQDi34Vf0QjL9F0gAV4LCCuC/uBXc+7hslZSTJyh/+ZhxPEqcFH8
NpSOFNXL3R1fdgz3pDcRN7yeqgf7nXZoWdav0cOYzxyDnDvl59ovWy79ifpAcpDIuIlgh7vuYjMx
//eHhml1zDhCXWQY1tkgXrqLy5D/5WXUxNuYKKI7x7pkPg9e1diLVVR+1rGT/QF/mcylVdLiLBB9
Y5yk5jnuYCNNYSFcip8G6AB14I+EHra5SsG2icEIRpSD3gC+wLsH+Och4wcQKFLnflHpLxhPSiI/
i62a9Do7FRTunC2ZI79GTZiaUIntc4Hev7+kMQn9fi7d8pI/2+3nRRPN1bCB+8+9CK7wVBsO9bqy
jGz7ZUnM+Y09KyEfz5h5tC1V269A9bires8FzRH6nYQTSZcKu6rqWTaVv3uqBrZ/tfAt9o1ceYIN
V6Ff+UiVF+ejWYJL2qZdlpSCI2Xh2Em/Xay/FlnRi++d6GGvMgqZWiMOCpABDCm60Q0uh3rA3YKM
3Rq63Hf9XTToUmm65MAXq0dtTh3EvbqyFLZ8BjNwbjR4VlfM8O4B6WwPZNFwI5PPb/jPMds8BC0r
ro3/3wfw1Jg75ZvHKFQ7F1w5W3oy/F4WC0XK6PhDjHvYVZ2iyPQPRxcvUqS4CRNIcvf7EcJcYIjU
Wgx8i4xbg7EbjL2Sq7wFwgS7NzgQcyBVZPJ4hXC10gfWwUiTYHj37Qc1m3JYf64lP6Jvyc0sMm6J
UDduT4tZhRs75N8LfawFNYcMJinKMRyxIp+qJkChXs8Ux/EeRRA0jjKALGOzYfefznMc8sOw+aqK
SL/XybsfNCDaOrbNuCG1M9XuLSIt06LRCUKb4uVVHMDkt/x0/9Dri5nhZec4Jj6Vrefufz/QZeM7
3XxH0ex0wfVGRysprZvpKmSgj25pkIBCZ43/qfkZAIYXyfSU0mYgOzgYu58WHMGAYvlkknd1Zm18
GZ/y0YpFydUWxMorDiTZS/+h3povazx2xVm8mrs3jsxCKOOWlQ44Wcv/FvrZUZT0DjNj4QIHiqbt
pGTMUgmYsycoY4em0O5BPe4r3cnvZIYYObLidrN/Y20IfjrW0NFYKIYaZnQs7KsSsM2wsMMtf+9j
37Er+RXcW5gW3zsjPfVv0mCOPN7xzaD2TSNJYLOmEgwNmJOsKoePGRgModg7zMnr4KxKBJfqlFWY
+0R3mRt+GcWh4ES+7kapzk0Ff5PgBt5PUC41vP5o/sL7Mlz62BwLMr7qNm7+bfsTC/Uv7ReZnbbi
HMbhrd2ZWGRnZqW1G5fzAALVmunUJ1F6uw16gE5lktoY8kVXsisu0SRSCQzB0RFIxUoVNx+ft3lZ
FoBVwRGiI000t5pLghpOZWazcOZTRi7u823sPmnfmeFZGb1p8fSZzeYvqFFNr5zTHlyu4SUCSez0
B1kg1yG/zdZANIIQyz+f+GVdfvzZm3bwtut1b2zKA0KG5ABrSUDrKqATSBjJribSkO+1iEOuoGot
nR21WJonr6LqCxVxCksir5F5guW0lZHDJDHdhL+TD3J1xy1GFnhmnRxfEU//TNwx68I1omBPvGD9
fNq2tRxtAhihB0a4Df5mkE5Q4tAHo44BppQjnK+gpsQfDDk2rBKjdcIoM33Bm+Px/GDDGF9VB5U2
kJ8SuuNsyEXkumKqqiNVyrMBekcSvBwLGMNdyrml6SmDguHOK5RPcoxUSjEueyvCTUrKjE2iD4hY
HxC1HiSsdp7bq3EsN2J7khOyfdqqG+D4nBgNCL6n6YrzjmbAWPsllFm7KyNo7Y6Wqp6fnzIyNkC8
dD7aLRs7YRnir+Oz+hq4dGHEPDgsVTF38soEL6IADRMaaAkZBYRrplySAW5wNLr6oNtFwvBXuPn4
eNt0Qqnxl4ZrG3P+RtzBBMYDHp1I9iqBafjd3vBEcoAYwMZTJulPdMMK6MdZooGaj4PVVA6GJirC
GJ9bsYzxnyEYJCnCEzHYi9vCJtSaEGZ02yPm565iqMJkwAPJyq5qCH95L1TKvKtSB5GdBj/k8G5Z
loJNvNzF26KsAj6duYIwCWUAA2KTZj7w35kX9YNuEk8CmpiPgGmK8zpdu+tP/NJFSZTudnGKuF/r
xGqmRlhuaTNeZ0Uf+BRCx+sM1L4PtvKT54ZGLlQsPrCkiYZLVukzea8yCemfG+tzUv94YDdtolGF
PNkZbooedWQHRBuXw5dcf2v8yBW3VU4zDZzKPmYjyC/S0oaf4AUOT3UOV3IoIc5ZzRQRbDW4eqx5
4eu1zGuBmOG6SzvlZVSiEEyma48yc2uXPAULu3dj2jUZ6bX5NvKSZWgNGTEmHDmNVUokNPFyL2Rx
Ub4nVRf6Y3Jw2dsnmYAoITT4lx6OenZG6mtwsQNo6zczqcR6J+PohIWFaTXIKFz8Ur13xtpf6JOB
kRVK5CA1BGK26o8FdRFRtH+2jWb02+e5hdpp6BBT7scqXaoMJ/P5RM4LNEirk+7BCl1Izrr4NZ3u
xZo+3A4b4CBj4AXkcL6pieHhwgPOJS/MBU/EzMTKTmyoYDsRcexLAwtP9VP+s/JQdr8KV1nST2r6
pGI91u1XALIdpyYeyBMBQkX9hudFvibb9U/n9FQg+aiWDcFqsGNbFke6Qf8YD+7cCq7dberbzP8E
8Py1QCOhd4ZgS1ak1ZzK2Aex6RR6fXhDR6+OhkANgMIVRhbmNtQkVKktj/lt4esysKpyRP4yx8x6
/tW/3Wb9e/+1f3NnIrzC1AG8bCWm3FPuT7MjlG4i5fnS35Tcyy+ccof+/hWr8+spf1CpZaliwkm7
0TiIVhRRdvnbIOny5qrsMt+V9W5w0X1YtbTizjKkFitFLFuYBDWw7V0sx06ESjwx+8L3mhpqINno
QI87SNdDKMxTNlZj9sreX+XCMvjCu51HygluAT6ZUdku6GBKb04og2KuK9OUHnzrCiLuj73yB+zm
x0tZcYXYZy6BXJIXbJUx5B1bzjmxyuYXOcoent7NDtMWy1UAiUIUJjaOaYLfzGQLL/ykPDD8J+GH
popP6GZipW5dD+IP22vSesAAIu6SVaLwNLM5dbiy0TsfIhrxsNY5ZRPbemisVACYZpZzcp2iTo2F
ot3yBAAXFdY80i47ZiI+UC4bUtia86/OpmN0RqJdhcqz8Cul9QfVHD7wosgkRrY7DsjpzP3rf42I
9msETB9EGQSRTfaxrtIEYZxdqSyNjXkuR7DJtvD61wHtIsEOOT/t/5WqdgIiU/k1LFf213YBJ4r+
jByMU86MLNPiYJ77JoODeGooyZ8Ilwi6vWBhEmmPseuiQVqgZcWplKWXTzGo61H+49pLFs9YZLXT
7rcYy4p1UeCHuzqaaKqZ9WLnqK6fBsQpDJQ/85UrW3TpYKrb35tS/F3J8HX9pt9PwUEvWcc8+0aB
8lvvFprw8LdQyZ4RpuojUYeHq3v21LNHnatvwmWGO564gu7O1VwCbHplBchYBo8Nfxg12sH9tMs2
HD3cOeJOFfSI6Vlwf1mWepjtmWtnPKJfO6/QQnxte7zbq4U5Jqm1hcZYyF1m249gc3F3agQFQlFY
EiLywpNb3Q+AESwP9m0ktRFpoX2jojvXEWw6zx7Kfdrvnqg0nOHP8cNL+4YsAdbadynlU5LHT0OD
l/mAM0ggDwlnGOAkF8mYF8cKPw8g4qocAqRRWjOqMMxGBIGvFUMMQ/QkV4yfcOrRO62KbVxmq7Lz
ncBtCgI13VXijLfY5pzPPyCdSMfH0LN0vyXBvj4C2Vo/0lApZYa8jR9GXgT622VSPFgaEG/66Z2S
rdr9QzpSqboNpAIGzFCP1y+5Lm3r3ZEP8PJSlnKelyTuAKTHxe6NPG2gBX3i/XCzlomORK2MYzUX
jUU86TULjmH6MKvlMJMU7w3vsrLtPzEjrcG0PzJExEShxwrvfx2PzkBFcYRRmXFRuaGInCyzoEnC
D7jwwqYUoWB5XdjEFAoRYVyFKXRhQx7EqgVGs8xjQPLMgzp13KuSSSqH9e/fLwXGp86/c4itXbm0
OGe8tY8xUI6da7TaUj3wcOg8fFTziKFuF+SdECYfDsHq61tlzUvlMDueRG3CwutWIl+35Mw7a8hK
W/hpBQDFaNkZV7CAS9AUeOYGSWQ9LvAe9qHtWO7UJELjksl4xtuyv9dfSOxpuTVYPxzsRS+vLON3
kthCmgmrZmE9n0KA3IXRW2+OfvSJfhmaBEl+5eOBlVy4qtk0xLBrftF1fw66+huMi3VjV2sxKde8
gAWBAWS6NpOslDZwXw6eo7yoA8m06a9fj4lC4PBlx5SRoW1QLeApbKtjop/ro8kKxkyanhzB1LJx
kV0VEDuwJfOkWAGyuc24js3YdN7g8Bqd0yMeOJlalztB34HJTa4Q3WxHUnAkFYK7htkLAL8dFApS
nC2PQUWaqVwQsEkBDWXoujvkYKhVASGoenNMdcHIMbegBWd/8zp9+BmHK2RWOTl4teKpzA961P9T
TgcGNs5TyM+F38oYhAXV/DrG+OOBbaQ2Q23e70Y99T9d42xIJkDVjOOMvZ2NRi3sztaEemRk+5d0
a8lMLIronFWW6SL3JQ5YE35sCmHoxbXPCyfVHv76VMfPvWMpIRO7ro2ZRQfn9hrtAaJnMN1TJ7tl
rAAf8zAFjCdgaCzEFXt6XtME0pc/yDaiEzKQ1ML/H0AfH8y/zt8hiucTvU7WyGUyxiNkqYK062zA
gzm3E2iMBFbzUrmNr7LQ4KwP5xNxOs6/I3Q30yPllLU/k3ErJSlh6Nm+n9Rfl4iw8lCdILdOfB5c
DXDL4yAdXQH5q9tNyHz1BY4hAL1zJqM9iPFAymL8NgT8vVtuozKFsc7eG6O76HF0Y6Zf2AgVJBMU
T/QrXOr4FnNr6HbIlbSrLkNotZLeqMAImVLMcuR4UzL+FwnxUsBfoK5LBv1Vwqv6tDXZFS2Lox8J
N5tvQ75br6J47Z/79mAS2psb9d6BATpFD7Uo6yrKseQQ+rNUVWllj7LgmslLZx8HSdYo2vsvrW0V
uWiyduOlkj5JmQaG3PfMPeawgSLs6DQf1glj5wdTkyrEi/vziXqqKppmm9ebnS+PNG6hGBY8lacS
On+DVFNGR8F8jbRU1nGpvAEqVumSZUIne/1tD3PeXbM4bDXEwnBtKt57MxVdIWJYzWeLj1kXARZv
rRcouLCLlBuUf6D8bUoGSQcAZvkaWzsjeDbxOQW1K41BMmJ4HrDI9MNHkUyvrQ86vDTgiFdOM4Oa
8P71BzBn2/a2kpF8AcAri0Qn0zMrq3JKcA1nLOH8iEpVqIFlVC9IY6Sgh61ImmaUSw2QOut1F5KC
g5zdGqCJp/eqlxkjvm7ExQmSr4Jmz+LkWPftCZawVBlCGqTYGcPRWKF9So4N2igwXXeF4bKSl2bq
H0cNF7/9oxOe4e4JfKM8Of87p18/VTKN/9oHIXMT//eCne1iljk9XNajb3G0n8tqrAokos15nm1l
uD3jaA8rQuzp/zq9snI9n//zHRUrMELzxbEnL5hl31Jz+g3XJT1bYHONaxAu+8OtGphJYPmfSjTk
4abq9JcKFQDvwo2Tu//EMQoKj66PpVzfRB7HDD+BT8Ksr/FrrWFi5kddk3o//4+n35Rt8DQ6femv
jyfUNczlyx7t6vvV0M/pyc87MyHnp9FfJ/GVSfgUT37y58TUR4hzjRb9/mpPDSYMRkuOwCeBaGPi
3IlZmwP9rtBRFso04JIJ0ULUOIUVj+UToRQoe3fQHqz/+HRlBZDGI3jvX5Ieq4Xq7kvsGE06k/8P
lCImI1KOFwo8vv95yzmiUqNDvH2H8EVZzA79vLA7Vqp15iwMOPivBB3p9YhJp18Yx4RY8DgiUpkO
VsXIul33EamX9056ceVdjoBBEo67ncpOzdjaxkpoHG+CEvJ4hKdViZUTRvQIpEw0CuKBfqQT3Cx+
TFdGcA/RbHR5DWobpZgJVNy+FyaknRO28g/awLdctY3FK6kA5N0vgNMe74QDdC+jrjr0AZl5FnAs
83TWoH+GbKzWt8vP1rXZDj5yB5q7Vunnka3skcTKgRmD9S1pak9oSlJMEJKlLsLPIFuMe+2H6QL+
6ABLd9gVTnHVAEkABiwMskjAjLTHWsQCn8oJHz3HQ4QcK1btY8Yxs0HQhwYOjyesJYHhySc0aJ6z
Zdy7liEJ+uPIPBmEWIlhvomCo9JnYH8nFF8icSmlxiKUljOrdocrNQ2aJ/DiFSKzuu6NPK7nsDiT
zgUoW7z43SEb+114BOqKn6/Gfb2/VpRuaxau3d8JjTmQCr70kOYs0/GSP2qIZQ//4J+tLzFCih1c
pv52tBQQehr7AoDSryEIGoYqAvp1df99VIzNIGw/p2gbMQzIY4hA/VwuaFy8L6bCyh//Kk9BSh08
quEHvQizL2mRcMERbvC/FeeS1vyKD3H0r22Rd4HDM8p02sMF27fkhpCrfHvbOMxKWlZ5Yi0F5BwG
YjU0813abAicWNUDS0NR5U4vojMfdFlA5oclfuQjs4vnJXsaYXBkYM+clz50vRSZ5o8Q/Oql5FIC
yPlxNfLf/oY5WyJt1GqSnh0xZziiZ1uh/0pIbnw/ak425mC1kouSYacvNDbewcF0mDimZNePOHBf
iURLVbrs0q3HObc7ipDslHyRyicQBMUx7P6xcNuKRZK5puTY/BE0sr33vgNt4TixUpzpeEX/t34V
cwLyZibLiQy3WFTxAIkYIiDzV3VZz/rw5ZHZYZJttVQUCQ1mZujeZUjQWrW1OD1E9YP8tKFqk/dK
InQzTmeifPfzQAL/dsO2g8tjKsFIPX7O/Ku8gWdqKdCNH8qtuy/9EuakPXzBBZxBQPd4+BQeft1m
TK7/TDTk8EE1FhPEhzsnqEUFWF+7Oc/xG02/aGSUXjXXs3xsHbtlySWmLd7YBqJbUZ+yIvDo6Wh6
S8upNyjTkdk87JKv+f99+pEpOks2pMl7/FITI+22f98AnmAIWbwitthBYYdQneBxv8us6hsdPRrc
m2/Mx1CnFidZI8/crrzpIIBx7mD4ypAu8PhMSPArZNhxbNLk1avYwG5GOEuvYkzTxM7CjBIaJ8vW
31GHh40KqzdudWxyBU3tnnoB13OxYh21TTOcEYn1FxhgvGmtJ6GHHAPUO4fTwt6C9Kzo+TmBUBul
y6o1xAZYeg79wKaj54FeEyNMYXw+CLO15SDYC8hSGQHyyHwClfwA9o2gJK28a1Buh8zu7yiE3Ihq
0D6QiouvQtumGgB1S6xBQ+TDGLvfieWYVln6pH5haZKofbiuezMDPLfbZ04B/QvwPaBj2h5kUeiS
qhxeBpqOlCN8KBgBERZIuk9ORsiWtFPXm1JJ08D2kebXFZAnheF3H6C2gzo+sTt1wizujSbtyZnR
YoyWFo2kw4/N+D9u46bG5+oOEZIELBMaCBOgCOG2aSFy0585AQXKDBmqpdMGjUTK+QUjeDnwAI64
FPFu/32ghJ6Hhfj/6PuR2SMnaHFBxkgU9LbfCueRI+R73DkYBv92jcYrOuV3Cxbp4E5x9x+7DNqC
+NrR4er4trarJzfe/Tv1rTgHlPfE0fFzo4Nf2rDSgF/sW4xgyrEzrO/X3/AeBZNnBtzZkJ9n9bDO
aQdRxAiv1NQZejzRQAfoEB6qrGrqND+wuvXox0c+2ZQkBt8PiVIVdy8HYccvYOX8UHtXMBUYZIsw
bGC4bJcPv+fQp5TLs0gagvb4c9RkzJ/YscBi/y+IBuMFzt1vS3eTag0Cax0j9GmvDdIrSchkL5w/
SNEcSzFmIlH6wPPfeAIPrkCvuX9zxn63Th48hm3ly7C0ab3/z5IC0FhUByyH96O4oX1uVzzq+b1U
LfKDLAGOy1JY9UlunxMnN4uB0T4RPSvgkgUHpfEV70rGLrs+pmKHAB8viJ47KIkS9Dq+62jsX0tK
pcWm4z2s/f50ltFotweqmp6K8JviPkoQ5EpzIMPOHspd7/ehUhfmc/g7f3puZQX+pQyqzFhJaeZa
bzTdSyrfgJ8eTPthmmkVCeb1bMSTqYXsC2pMegdrpnau2Vz722gMsxpic56iub5yG2JSed9gcyGG
BQdon7/6GCZS0m1GZ6SwCtW6ars4fA2z4sm+roL2GeXiL4wppCEk0a8D9Ew09plBytyiDvVZUCLo
erJKG8Tk8NodeY2Q7q+FXr5NVcdzBUXXfibB6x61bX5nsRJmSduTUTuXg5pbTLs4Cu7WYrDkYCYH
2nSfVhVzTwLqdCg4FtqIaLIqtTuGJkGbZoGSTWoA1Nvkd9sxf4GICS9aWyKWoiGj8Nvi0Q1roQtV
9khmhOvc90zLs4Q5rIPwT/WBkcs5bbCfIsHcfD9Dx54rhKiRYNa3TRgL7T+xoqbhpX21at4odh1o
EBH4Dd8G1wuBQG8kmRFX1D0UOHCu3tCgpkyXduWe+jZ+XrWP5C5/yd+vjqed+unzf6D539y68QCw
pqF3asw5z9oDJCbIvKDrm2b2c95L2VkAkUy7FITqKYWmsHzMvN8J7Y02MfqK7sNkiib7wvfsm+VV
M5jTWMV2yvpbcNT7mcJ9Fk/K2S43J469JYp+aXqhrwdB0pdlNB55rAA4P+5GfUlu2Rnf5gH2DT2S
zoKud2Q21LKWW0uo/jsjq0IbDVo0bn6DWey4bvzD+eQvmpwtLF9YHtJ3507mNcGrthFrEsa16ILQ
07fGqskHZR0aa33MDfYUOZtmxudsd+o2zAobm/WWhRiIfdUxKX5N4Ac5GIhDcoGZ9hhhOlfJE4wh
cRq2mjESJzNrG4OLAtfzHgecTpW8g1nIlTXsjgSp6bbf/Dc78h1OE2soE6XNLJ9zYOReyIjkHaGz
aYLmNIc8/rMBBIoQm5ADNcjvZ4wsE1WNvldx8Q5Foo2InjVsDO83wEezNPn9UvhmZEYT1Hr+/az5
qzsaZCQIB6vqmBmQaYAHiqNslSQxmVkk9qbry08ZJv55FrQhPrCTN7yFKrZpRQrqFsPjhPKVoBnR
V3FjQfF+UjUr0ulH+XMOiRM3mddd7/Pg1hEeD/aLqiGB6pa7eIqCVky0DI53+h993t28+jLkdN9h
m7GZJvwLXbKszNlz7haCHiudRVW9cclNSA5kQlVrEjsN8b03sbBHrzfPvZP5x3Tg7ysd2N+vi0Wv
fx5fj9h6lbX51p3s0j1gd/GBcvUu4SihwPL7+kPzvRb1afHqMSWfDn9VFbB/Kd04Tc7GxW6e0vo6
jSaBamKIZ56Y4y4y4EFmBk6CilWAOUm1ULgQt+22PCqj0RL+OS/JRuIpeWvaO69coutp5dBEHJjN
SwXzXaCZNYNd4PpVxmRBL/rXTpyQRJ5Ij8gdA5N5YXZYIrXk5nH0g7abfu2F1pvuL8rqFG/FhBzv
kOqB1Xua8jMvqYAJM4PpTLg1OkzItyETvWQvuzyNXqN77CpqPQuuXMYORn+oJPZ0tXqH5umy7PXO
4vhWohpNWCm7/G7JlMBL3qT7M2kKCkmskh1vYqJNVx5sFOkcmKzx4LuYSsHFdrmOR5tdKOzRXGqh
lQs7rmPMsvhs59jB19XvculbHqRdqATU369/UOJJTQtHOqXVr/YrprNghQE7aWeUspQz6cQGtI+H
mOKLrlyoBENzv9KDI6VjXxHARZ8Ech8zzq54m5kBjnb/8YBNEK+yC264vFhTiNxLwDDdrNex+Xlv
k0Tvn+vD51a1ZLQ6UbheWlo2mT9IdqSpqrpVC5WSjVRsYwYSxTl52l9hiTEGM66dUuWWB8pY2vwz
gExfp3DIt+l3+CEcUirEuMywf2sP7eVn/IyUtZlGpmeBcjM5xiGuGb8+vyYD/s1LKqQF3BE/eU0A
aa8RbC6pUII5u871EcQVlm9ewFXsBM4PEQDifMXNjp9IMy7f4Zn13luIccwilw8ldQ050CIpa3ly
5y1rAub4VDw0BK0aNfDZX0h3InLlQnQbkQtQSx877V923BBcb6UGHrK4w1EAYtqj7j0tJxiWyIki
pvN18tCPFMOrS24HHUP6pYuLQg06pqeH3FFYdPoMC9ejixPJQEe7wGvoxYwtKh23KPI5xBoSg1Xm
y3Qq6iAAFMhl6R8h5HOP1GxNOlPvdHQRP4v8NvYgzxHuQ/RtqtjOXz4RKWas3mGIkNmqZcJFmPW8
wCHYwAXORRn6Iqwc8cmmP8LivypEbCOcAMCAN2jPlLv1dgjd9BvmCKqCCdkTjEY6iOsHIY4WSENz
/dVVcQzxe1cdxaDHpH48ZIP/TjisF2TxWq3r1s5CwOpglNDqxvWQxxzjBbyztTl2PEecY1QOeysU
ZH9R3mrbNitT0InLXEuJjM48KN9/8uepKc26w78EhPa//tQP+21BhRMqOIcYGV/Ov7rmjZZU6AwV
rwNRwXTPebQFUXzSuUKXUly1ga577LhxKPMBVBRMnYg3W/m/xDSEKtFpV3gGYNk/gFCHBKYW5g2i
JIcEYNwoGMoOAK72QkSoi0xeaJX6xXciF/lh3Ac7LAUz+3DRohQRFvQoxCaEQllkMsNjg85JhAOC
DC47A3M7vHfLhamnRcBmC4MgHpCRzmDfI8/bmEoWxQ6AJ5sMRKCI5NBSi7n6e8qYrgDupeGMiXwg
ykpyO24s4AbyxovXSolrRs13wWGxmP5yyuQNVy5yAu2OseuZcR64/Ymf8BaTOWlE8qFp4J3Modlq
LqxOGglCalNmqPpF+zFpBbem9HqzH/KrC2bcgofWkoXIWCwOVoL21iEKdeI0mOAkmTBk2rTJ//+3
TeZ1i1UUDRbDcEQtCGgsJ9n0xsHlI7MNn7w5oIaXN9Fjz3f33PY8bB2r+LBDXboaeixd4ZTpA84Z
pvkEy1ayQPh7MymKfWT5LxLOBnaJR1QSo6JccfvZvDiwHIUK5skX44O2oHAtysrNOXfM1MC2B058
hOpJvmbNkzCaf7O1gZHfZDLe70LSJRUVPYn1eTwnyqJnlxeREDgYt0AWENDbFDJtriOgRkERqmw4
dz2JKJj2lZsEFk6PCJ0/pv21MSjd/WBz2N6tuAyvEm/lUtQ5b78yXuuoCVnerL2zOzXp9fWB75bd
LQkNCJ9wztjGsJOEfG9+F2EdOep2AvSMT2H81OQW7fpms96WdP85/0wUnbX1Q1MB+183ggnUi8+E
IyGwdJCjO+kt1y312oqUiLiiiS1KOhS4EbSgj2nQI6tywa8ce2pfvSWj6197R5iwakrSAIF+xWyM
gLlsiFkkvuSrq22MmYBE8Q2frBzchyq/EAaPMBJ/6c6VHG6gw7NXGzfZtKqhSvpzjJX43NoLq6l9
m5SNFGPvBv2MAyy3S39wQNkIgtxquGIEv5aUvf1VSukRjJG2+zR2OXJlcC/ADsNron1JhJnLoP3X
3lqh7uKUA+kMBRofaRXN6vOSHsrnx2VPXC/QGF1o6yQPPlrrkBuMTEVi+8TcZ/UUMlLtF3JySXyl
8a2zsohyL/04wgD8PFg0ItTl5fTDt6F5HdWfU9YiGsC0/YoJkTR4Qno4Hn4wxxsSz4xJLDPxMaRk
hYZTOWLP4jFFd7TPCeXlM2Wl85anNruPm40clwqlH6t0bjSLu+LodoWImrOWhK6SyAIh3ZJJDO78
6HADKgyUm+MO/V83ahBs0oerbZQqG0GHk3bzl7wYjH0Ft9wCtOBmFgPK4OTkNA7ngOOaPHH4DZrU
qhNIrsCYgT5oFGH84Ao/imYvP35NpWuuAL2B6KW+dJNbtRoI8tereg2LtryqQbt9BbJq8MI9rqe4
cIDX3yj30TST+V5zasYhiceEoezl3rVmGV7WhdevZO8yi3bXYgV77nFFzkLXc3/qKbd43fexLKqu
tRWWv8XiJL5NdK4c5/qbRsRQke8O6aVC/dgYrKsPwJhGp4R/gsyZZYJGEpbZyueVxaw/lE6trcan
qYe+wn+swryNI1Xgk4LC3wkj3eCDTQfkA8afb8sRvXe8/+SXxPELsCMNiCm8Bg9eXQCl66wV9Wux
5VIO8LzygiqZd8FxLwO0TjfRAFJjKj0vAGqLnIi2kGnMaIk75WSbl7PO7KiHr4rNlJQeXbI/69zr
I6B9AMDFnJVXTUCd8JlD8O5JJHKmHpPW5zAv6BT2PJvtmuIgjSCqbL0B8oXtv+LKkOETaK3nKR5u
lGbUj+PcwuYapohVawnZsuc/xAdqeCdU1Ef54z1FbAu4TCNP98zt4FwueZiz65SfnbdC7w1Yk0gz
UuT45lfsWVPoMghcCzfNx6FiSZhconMpxwkTQHMYdQr+aZMpt8w5CFa8drQmunnxGCR45hhfD50e
5Bj5ehjr/NEYMJ5x+Up8Uk/w7hgE6rXj0DP/k8m2puvcCmWB4ewECYHWJts2hfs/ZhCX6ELtnias
4Db5r4mtzemQ1qSjoQfrqcoljc9LFeuD/7Wz2wQaX6iTGgSTGzGsHltFWBGqVqIwONKR6DquX1GW
3ZpuiAXP5jU8YpQAPvVDD6rBbGWHSq/R9XJVE09RfvNhflYLLTnquWRCdR0q8ygd85LIiUFEW3OD
dRCLO0ClDpI09ioEc0qfJfEwEscWrysXnXzTBUFwQxCrkXsJ+sFoc/Nt6w6zCLcbJqLmOZ/XvQo7
uNfklibM4AtFcd4AJdHmxN4m6M3m3F2hpk5jGQ2YMYTRrs3ibk3OaIp6IA3IGfrLEOEsrhPhZ6NV
e2GgO/XfxCyQmggfmGEoEQL08GBHgAb7Q66n4AN0KXdFHv2EM2kClQGK04+XOmh2rZz+FHo0kFJs
m5OgKhyvwI0tnSH++Lr4eoYrRMByTcGcetU0srtMtJ0gDFZZW2ur9WT3zPPTaxZkpZ/EhAXNbgDK
2LASRqNQ9km9aw3HdWIvJggu3U2xJqOkpdsvEZQ4MLCa07SxT4NXa1Qc1Jkk56qUkyOYnXKbCT1r
2/BBKcaa6FJ9af76uVkxD2aVeZzNR/76QrOo04sQppa0cuSKLHmRsM13LKQevBJx+6Vj49/D80D9
1gkWubwE9brk9TQ8ufVdwbhXQwf6PX2Ct2e/lLAOVKuAnOcdLOeKYPKvxjCpMPL4fXJ7cdBGF3ol
T0o2PCY+GA7MwrY9u034e5xb1eX/VhL99umpDFSYiJpNiMdff1EW98UxANpkx4K3KVtd36tb0pqc
2FXHT8II2uahGeYKXLMvC9P5aSv7fbxE9XpXAHd3WUXYnOPfCAqMJu4wYaLAMmx8fqBQBKOr8YeG
9CvYd9ko5EGj+nAWeC7c5jZ4gwc7ZjERdSItlrvZYfWJ2t2B15OUcvjcpY6l4B7NnK+SsCEelbEp
4lRUEMXPM2qxofHVmaEGwe3LR9twgeB4hlRZ5FBjyz51Y5CykoKda2MBWrnXvEqFDXx8aR0R5Y1v
vnY9O+7ufiWPX4zyZXp43VHlRMWu3DGxHXYlacMHOzTG1lbD9EYhkvUzG83LFVlYzr3pBVf9bPYW
JE3qqaWhxh8tXROjL15aUT/QqSwuvTKkf9g/6+MBCL5NYmmSwv3AnE8GTGJiCHZq3BZW7YvJnMP3
FeyFDoEmLRhWUX6iJp4Q4Yb3fdHjGfTq0y/AnmHJk0QmSLahQG0qFxMTBhirGeMXAvh0CiKxvfGO
W6nHRdk1ckimz9P7y66u0WY+Xrhq0UgC2Se/WXgcnP8XKVgLBwIRrFVhECxYj5YbFMYXPUp0idc1
i/fk2njvSgEz/izmgI+v2m+fdUO4FAPgjRSsFpAfArai6tPvNeAde3umZl4fuuCdEnUb7IZ5I+Nb
aWc50PA7s/Syvcjj3crFDG6QQX1TXJN2I+kiO/XHYI6MaKTb1rkUKeDtl0dXKNGinxODYPW40Ddj
LAvC253invECxheIYLKtpr+u+WeTuyosoMyM+4To00eWre8hyXC8xvIl9VyAUTQG0qAfpQYFxGS+
0Mv0nGY+VO5kHF77WKid2aX9UKpHXbupvRUikvKpIRma55Zhb8CvNOlCLiVCuaL44/ALTfyW3USq
/xoPZMSxOZxAQCIR/V7seD9/LJaGIx2rPKXu21lJt8eJLQLp0rfXcH3m1iPstYvu6WJDnMi6Akt/
q/oZIVm4GVLmLYxYFBZ0l3CVv3j70FTdQ+iMJpeSKhL/dORDZF+mIl5QXxrd86oQlfl5cM/NKAl0
9E9Z3pS5u6o/iIdL4scCF82gepU3ZWd4GPBfs8zrccwlvrj6TwpQwZmDk0NIfSgDAkILw9zOBl76
+odtB9D15s+VGCbIBtSjbTM6dBDZrZerhZJp6IwtuaB1NcgSk/DOHC95YTanMgMrDobz1v8HhkFB
IB6KSj/K2nDJQlsmUQWVizlHo0SRPOdd0OrwopbgY+c/Tmd7c15d9yP1QXy/jn3fJuZjBBCZaG15
9moJ/U5d+Mb/KKKeZWUkShigpUXOEZAgV97/tE/w02VEH91Bzh2pXeNdjbv9U+ueEsYupzkbkWZy
BsIU1/k+YwhOVfDutfPThHBtk3bWY2lWohS/Ovi8yGQU1tN35EEUqzHlpktPj4ms8ODWgxpKqBO0
zj6+VUYgMB5WoTz4BDBKlzf1D4pa1J/49AydyHFoJ5nQ1GguQWO7fOTJBJd8WJRJwLs10TXVZpfc
inRVIuu4YJNvOnwClMKN0LZ6TaEVsvyncKisK9aMqWFY+jRgWKodb7sbZxKR96/SywGtTeIpP7Zs
WxRfTOWdTwhmQQr1lD8CPvZwRhfqIim2Z6bpNXMBSvgZ4I80EI0wExXITSsq++m8rVlJAm0ZVHbk
fwGHh/5/N9Arc5IDeRLLkmw6S0aysIzBPC/ufEOhVDIFsJXpnj03KPVmpQQLQOjhYLYjHkI4jeaC
v/L1tOfh4USQ6nUByA13XLnwLaR983p92iV1w3dGpURJmV8rPgbg0MPtQWOtYljcVhxsFy8av1GW
mYf6KXMgZwiS67Bqy5rNZIeK0VB0wgZ4hdgOZ7ji/r9V49J5p8I+LOKB1Bv/yKFqPF/PTp0FYF9X
nLQStAHsJBDASLtT0wyocvZTYOGB637kpYPX2ptSdmUsTc2XzTtuANN6GOz3+l26keAly8fg/hdY
39CfIYZI2RVSYIHi459/A8T5HkfZAnjN1USOg8Cop2/Fx6NoRaiS2Zu3aInr6sldF4OLm3HsIjlp
Cywn2ujw5T11sDOEbf9idfG3MVng1CTYrhwOVWZxNshFm4KbrcAKtydeqnnsvPbLfQ/kGND9VRNd
+zPHmiZ3Avo/30FTUSL4xQX+IgoAtd+TyFr53UJeZ8u1fOQIi5nNEUA3J71LQ+j9DAcOzyZYtu1t
Nsq2EswJmGRF/r5heNmxFhlvIRdOk50y2vT29Nxzyal05U6azVGhXdZzOCBazF+0e299OmD/plbU
pFsoB4iBAWvOy3Wm/sGAASrPz6AE+RX8VNf53IJtN9va+cpA5hZzZ8O6CPyhK2DNXteiyuu7dawG
AReEpph7BdUHapLDkKNoTcY+Cj2BqQzrDGI+5fEHHfeyYHA1v48MQXNqmSFHfKhXMY2xmEl2J3bD
Y8KEC6fa1pIOjtHIGVimejLiSpIE7YGRKhsivL4fTFsMvD3GBTYd66YcVjXNNpG6iG/kauHKF0kO
hJSJeCtKBO26/MdFXHcUmBW2nsh154ss/tALB3QtiztU47Y7dAAnufsD7aQFmEc9ZNCYcqd5j3Au
DKkYWmTDrPdFhFr8lq5/1pOSdSg1lKX6cPQW0g0hCh3KPVt2tk/PL5Q9TjwjrOlPquINm4CMaemC
8Z87haMSceFNaM9rG1mqNm8wZo+LKoS97Ox0FVhR2JhSOTD+37k+cmp7p6YR33+bdEyyr3GdMCVw
wqCMJIgFxT/4d33D9K50BPAG8Nxq2Tuno9fxUGrP7RxV44uchyLKzQwe4EZQB/QOSUaJ6qbRyvEJ
sWTySb42KnahYf2hHNbmW6eQVtH5pYbj8ThGulqVZVdpp+77/Po05onGtanuObT4ZhRZZEAlsOrE
0IDa4KWjfFJRBeafTLdzJ1kqUIX7pJlbmSpU+M3+3OpwP9JLxXCIAo88nfPWr0x4blVh/y1qj0WJ
TtMqjVmWyHJUVnpFXJZAKZdyRUTEu5VbZ8PZTaAHXPpKNU1FcUrRRZ05mMVsJ73I4LbALNf4diTm
45HjfOlKAJdnx3EynRQvtXzD+NAm16Ifs08VulY+/gpDPLmkUt8KIEPrRQ8n58a9qonlUOdf6xt7
GBjDpmF6zTGQoL0aDiJTcjRV6a1AVJ617+XlLlOtjmrYURGbwlz6E6WotCOlku0D2G5Nsz4KiQwy
9JCECcdAziY/MOpn
`protect end_protected
