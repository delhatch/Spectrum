-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DEe9m2CnQ0L1hKhQM6ChKUJl9QVJ0+QiJYJZITHvQa23T8+R4iUf/7R/MoalMKQKXrbnBRCEjqB1
6EV5oqOiksO3uh6jimqgBmhcBFy79hZO4kbMG5RLSZfa8zDV1p9hgSjQo/Tl9pYaXvI3uwAYthAs
AJTIzjOoAQx552y024Fgo2tTJHEmAA+wc/4iLXymO+HVSeInmCiH54Ghsp3bVXK/vB9Uv5ZNMXls
PdbCZg/2WVH2d+vzMkMcWvBnvt0ujTr03mUbmx83XzRKYYcNeOezXxEd2TSeLfO+XBHsHfpeWMAA
JGP+zU02qb9uRO9GDFBGxLkJZmjcJQ7fUzAAuQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
fjtRkaGny+xHb5JObFA8j3m8KvVXKi77Wrg+5/m/j8atzzh/MDbSsxFUSgGnkfqkahycK7kvRYRd
UVOwAiAUaKuX7OH6imjlSVBVDvQ8zqhIyocMkYCDObdZFOc0HoJz98GPs4CpQGkvKX+s7uJ6vEfv
7rQQlFRrRnxCEXCtzrB0utcmhtVQ/78HeYoI5Fnwo69f8k8GPprdyz32+0UVKJI41Nkba+ENqsMA
8w8awYVFutIDeMFSSqrfrUK73AtbRWPjY9pl/b7krctNRy80nHmTAsM0eMpTeBGzYiG7lWBV7Xuh
i1GK3I9g9fE+TfnM06MERbsd71IPZ86fmmJYFahZ6QQUiUj6dwVVCT78aIh9P/L9WD7M/XDKAPXW
XEvFu1gokJTCYpAR+rJE9vR3jIBLEDeradScWRpFNClXlm4K77xUcIWNi0xIlZJcZlXTIq78tw92
MmumnlqvN4/gEByumEqqxoEfiRyT908joJxzvlLy7S/47wHiO0e575yHAV89B5+aon2Zq/9bWUtp
qOWJ/A6O2x2Mz2kyqfH3a4mOakF7SVKb7skjouZUdjYFA9NOjS5VBzX4VktIqYglOzNlfDCuqC79
0SxCWEKCFhVdDtdBz1xPThWJPk+WxgbZwhbBj5AJRK0AEZOrLoi5SQdOpE7tE8r06vSXDzB/5Opj
CGq2TjDt7jMsrY2Dy/Q5U/STnb9avnGjFa8b5I6E0mbgpc/VHK1+mwWizKp2ycXy943jruaBNBGi
hocutQMdvqSvDiDzsCUvlAkvTIynEJGxirJo/Ra0rcPHFeM74CLopUA6CMMIJBb0hR+3SxRRbmxC
jnWFofIZpb1tH+PB41UdrADIS5pAdIAmr8mBTvyZI+Bn2TanXJgJYR4tLsmpUnJEdDFo44kOe+kD
J+bwS46JI675TqC/5Aj4eQ/SMVUwRPd83P0+vEHU2CKQoM8FZ+Pm5JwuUyaPyIe9IwjlLdo+TKOH
vqwtW6TF4YTwa8lD2QTjjORzmV/LfnYdej1nzFBHKTA/q7qNUWVMKeh89x4p3r5HrKzFFKyEoLe1
dZ7+CiUiAu8vMlMlU8QWuoVp1bwnueQ1dgC+N3/JRga8wZrPX+b7BLxqKfTvPiNkNl01YQgdy36n
B075bW1FBTMIomfb86R16GN8uyrLoeZf1xrlW0aPig9gUDgpHu5owp84PIJyLrtCoseW8Kyplc2j
vrMDhw2yUSQATJzXXkE87uSJE/tSAsl0lSf8cCIGOr4kA3nARtqKYM5ksBauh3DO9Ysm8VVkJKO/
lRMaAk0o7vLMI84cPJ4SXWWXvHhAD4gXDihbP4WG35ipSLGHLFqdzKd5dLcRdCBhMzWq1Q7UqD9Q
o52g29w2QlEs/eCVBbg/KL0spr14HGvbUnY4EC1G1K8F0gwWn/pf54hIyg7A+EUkHWvdHA5MSft8
B9hS/1i/sLQAaVRKzgChHFdRe0eV9NNomvLH2AXkC2+IvteyP+Fgf4gaGLjOO6MkwMvkDPU0e6Sd
a7j7kX9YqER/yIWRGW0KhcuayjwcVOc1trzHxC0YU+80Knw75dGe8xLTDB8eZwWVkxhyHg8q4mxc
IuA0sqwfYwBSzoJKSlR9Eowai+cICPff3I+cKnEnmlkDrliEnFhY9lyfwPZR/AaRH+NcnSXboCkd
Oestx1WYCjoC1dZk3EtLRtnTdT+Qa9mNx50IOVNTbwdbSK36M2/WiT2ios3Ron49Koa8erK+SJAb
P6Sk5z3fsRCWhRaCRL0mbe+I7KPwFY/sK7exiWuwqjNkrUWi/nxfjsbWC/iVkPcLIGEnmG43jqQH
pDfo+askefVOkeLiTSWA3wErsRs02apuCH6kg0z147/ddYAj5gQXKYyRYZJTlO71EFKAjgCQ7XYU
ECan8fne2Zxvl7/dXTcQSl08+1t6aFinu5XrCTbPbecGmj++AeVIYY9V4h6xxrFcX7Ue89CurdEi
7blAM1XC9V6nRIcHk7q0vQp//fST3G5KaQFvDBRYR6JTxvO07OerIUQFzIek1+fuBSLrx62I2xSC
C9uKxIV93Ppn51gTTatqF8Ikz5MpSw6583esCoC2pl7U/P0HkO2Y2Zy0HSN6lH1Pdz3Ynm7eioiA
PJiNGIE3z0+PmQhlg3Dh+rwQnCemf6U2p9IZvTerSagCv98echiirNZc7JzMoPzvbVraJjNtMbAu
UySVnrpz2g7BUhmyRcGB4JboBS9AvU9sBwFtI1joZrWH+plQRikbKfpRRdO3MBSZG2fNvqVB9j1y
xxuQtvazvrP/gxeyK2SCQ1N2EGtnelLIQMmiwpZqhKhkdxSwGWdfP7lk0UIJNsyyBWTF0dPYUKxb
X4OyWhtqQzICVXWg70bs1O3eeG6FiKLDE2t6S/vs2MkqxBwSdgPJqss1RpaBJzdxUuWgLWpQElMO
FjmfGJkIh7M1cpSrLvJ1lmZmOonFXJuJ9yDcwgxZgiM30w3o4WSz6DOwynCMhH7BZ6m6NYalTGCp
5KfCvsVAuMUlCUNj/Szra7+USPTphIi2zIXPCeeEC1iJoOk+qG62t7G6FiRD77MG2NFNTUpeJgTh
fBTFw1KunjNS+X0XaUrZ1PHIBB9Ww8MAoek2uKS3jYPBYDRb4YFYqU6dsudbLmGem6gttLyy4Sai
RUd5ssuSMHLAkSkIsN53yzCTbwd/jkEDnyX1RoFP80+WMc+4jT1/Crpfl4sJZ9dAkB6OZBjQGxiS
V7Li13/GTzOQiIgmAIPzCccdbSxvuSAyc7Wxo8un2QN69glYs512wiiGRybViK51jvmVT9dzc2HJ
fQYnrFqqaZr4BjUMmtzuDcGbxAhcw0XFZ90Nykb5QVWNIL8WgWoXyZO4bK+azvRdCP05H7wTNYuB
WLMykoCGlcYyctDNxCBq30cLAPmfnWpQvIhjuAS7t3VR7XV5CSFLNq8vNLq+JTAA/uxUGtwb1VvA
Q8T7Ak2yApwVlGvY88OHjvyWQB55B/+8yx4ni8O3QrPY7c38TTR4vkI/yhInk0CfAJUhn+l7Zy+O
15Zz3oagpkFjvIX/nY26u47adsPC5JeFXeArMvqtlHoEXFA1PzlOsXXELlplupD8b4aevAqoV4d/
2KywzmCCOgc63l/IXzcLsiosWDVHEpU1mvhBEofxq3jj6zpwpNWvOd15RBUoQW/mnyLx5TFPC7MT
+iGhYrXXNsr1I8YAh1T3kSYMvMEWRqaBd3OspQDhjNnO/y2iBUzBeWhLo57AvBbdMM7PVwQ8jNYJ
+GXr4JAM19D0+CzD0iieJ+RbUsSjmpAifpL/5l1WDKze/XejMKIDWRG3bF0i7IcWz7FpEKSFi0Be
yNnp9HUWCCpGnCysyZ/qhyhoygom431RREFJFvUIUsjzuJ5a2+ecazBcXlbhX+mWdOjIB4dlsK0z
THTxzaMITQ7ld+Ws9/LqQ+HIlp2BOy9l+bElTivNrAG1wCEelVzB79Nw3vtEFRIhBzk8xm/u6F+e
SQ8T7AAB1Bdgf9idbAjg1fye3+Nmt/CMG8SvXknsrh39vtzBgjfiRNpNoc1uKaG95UMVdRccV5uf
j6C048FqTSS+4vD+4rO2ku6Ha/5CNKB890HDzqMT/faQY+2jQJKmQnUBfXCDW96deDefzsO8uBu9
MipWqFbT3eI/vfByGgZn41n+E7miOHxOPAreYX7Ukw5mSL+lFZ82zN2ryiDF8ibNkjR5A8yrRY/K
5zIaDOvwkuUF6IMbPcLbcwLJV6XoSzOISSZSR7JjedCAindVPU7Pgzp6QX3Dv7jP7M57+7XokzNG
FOEKcmptB5dBoOCUeJ/f5lgu9hdUc466K/q0Rne0s8iG7zG0GfrlDG0DgABNnILjaqFUla8nBm3t
VR2e5mC/zoFVLJd+mJ2IRJ+bzLYfGCb16EmBh9De7aAVogj5wxf+T66fPHkOo8pBBxv7JwCnMQlF
IBbd6/ZY9weGVoyoLSpVVRZ4cjnhQex+o/PkRi+esjP60DvteQjq1CcwXQxxz6Tlhoghx+fHeLJt
rdQE32Wztbg02XcIBCAzLgak+MjKFDs/Zu/Ktvmj1ttXFQFqsk+S0u8weKyNauikA/ejWpM/sSs6
C4wREpx/h4kAn6IAn1u+/Dm/DdB4CbD61aYdnVwAvYW3nJ0u+oI4WsiyI9OpI1afGhpYvZij+8MY
ibeHRJKEntlW7AY5vEGXyFwRF9Rv3k/rFmV68TLvT3THCYPSWLK3r9oEFmpAIRHC+LU4JE+meBpE
4NxOepQecEyWdVvt0X2skWd7YwDEY7FdLhStURJr+xxTQrjwo5/zFbbQWm4XbJGQVsHZFyj+rcBh
i/okv1WrK43PmxQHwbl1S4eneD2dhuKlo4DGL1oS4actdvJUbPmI2GfCxXK8C6GsG23atF42nVeF
NkMs/Ny3JANGwzAHMBh7XtwqhAxv0RuWnP32KLWEkRTbXaxOGulUyXawSN5pNjM+US9Zv4sNcHrW
THQ77VEfWcxeQM2VHhXCLHvCh8cPaPJ/E7khjqIEyCkTjk2RaWedybJjyfLwTwlo0t42zNmGfqra
pt+eMzsm+UNE/J834uebvdJXYsaHUHPnmUU2lA5JeFNfTWqSPFfcNXEqyuUS9CB3UeJaL/6A6gXg
1Us4p8LXYfgX0QohNYDKRZuUKQaiOUgMy9H+Gwrli5mdp0UcjrNcQ34sS5n2A0JkSuPoyHQd92Mn
vFnoOKiVMCn5ij4EPPwzkRR4vRNMgMUpFlVwdcTvO/+ciR/CjsxNWi13KfR78xTOTdCVCJ23Dcz7
f2Fn5Pklu/Neq03L/laefGo7lu+hamzdHu92Dp9V6momaW8z5e3CxG4PVXpiRvdQmEbv5KqKZ1tl
KGdZ7+rNN/o9h7309JZmidNFVNrTrHoZCnWipYM0eK5nM0v4RXfpjrOiZwJtmNGodRTMTW6txSaL
UNJzk6NW16pXus4yXGgOeZVo0E+r3ri6cBaTS/vs9Zl9GogskwGFmzBQsdX3bnEY2WBJ4lfEZ3oo
4eqF5MwdiukxjQ/JnqsUpJZZXkIYv1PQpjH8E7VAX0Etnpii2/fAzlOrtZhw/4FkYK7by9a01/V+
afYradPhMLjfN1b5DQuwUqHP3a6vD3gxIuJGQH6H/kdfMz5DZQ+3adtZgh5GMJwzcvvylKEsUG+K
DWXBznsadTgni7lCCVvJn+WW2Wrjanjhyhnqfuw3ArhB6Gn9IlRmPCxctuF9Eg2cHoMxonZ5pW3E
gLgHnrHpSxAeRqIWVJUz/0J9FOjQ4HJguVSvkJF2iKjnCF3Jhgv6EAFRJ9qN0zZY3zejcgbmvGBq
ZsMDc3ftyG3REBvJRyw3Cp5MvbessFKrienRpnO12pAnzUqc6MrBYuoR9AVUsi1sTmUg5y84TIpW
HcxdsLSIXQeNjv89HvdKfGXuAwD3RGvutYyDcp+5ltLH58TlaW7UNtEXHq8ZOoUOTmk7aYxR5ohz
PPF/HNfwarXwzyrqX8EBNULM22h3rvdzsEvFFlaE+bNza1nXm0054lwOVk2XvQq2bhWzjJqQ10Vl
5d8CfbYhdE9phuo6tV6Sd0zQTuY6luHvZuUD9tzGvD7ds6Mz0Kkai7PyuGjrxjTLULWhwVbFT2Zz
p94xwd8iWmhD+I4sSddFLLTeD0sf2vbmu6Ghh7HdyPo2ejsLHgKcSUp5ibJTd3Jf7+6HMK7o2o2x
Zjd0rkksz3nt0REDRvzNSgaKgm/Jbn9em84H1cFXaAzS0fXXtzvqyM+4gTbjrc+BSoR9NiWbS6a8
TzZeI6KDQunpzdT7Zx+AJYHRs0C7KpPA2ZY0rAchZm8idoBNCe3PcNxG7bj8C2702B8bf7wz3ebP
q7qwKfeYAilzJUQu77StcPunD3z52JCLeDAccwQn9AaEEvP4qHHk0AwNSFPWIBdqQXSC0wDqF09z
MmcfTLUeqeYt+cxZKYf/n7ZVdH2EYGmJac60wYfndxHjy59w8BbQ0fHgehN3akf4ys3qDDh53GWl
D95JB924UgzOh8rQC+HOasnW0wN3nIcFBXl95CTK52xHW5OUL6NdGiynVeUAPS4wYDTvZ45w98Id
2g6mhL5a6YIJGIZL5TK4S6wvJfv4ck7FDqo7vfv8yA3yKbrJvHJf65tiAq3d9jFLdTfWM4yFfYiZ
Rh5I1ftJ1b27azv945TH0h1oij5T5XHeDlqpCeYdKe3LCVjlaxMWwwqPytjmsbabICdfEaGFwEbG
OSYvzPhYOaxDIq4LasGFBQ5DG5X4ZcQL2ogCP6dSRhEgVYWcgqawZvdiGhj7vLUouAAy4FZriEZc
h5heIS0D1sTOauFit/A+sWgLo2JzpOABR1HRulooaLPPa0TlpSFTmPTzC8nWBPAkV6iVC5xZ9WMU
IW3v4jfZ6A4w0LA1lrFCj5oQ3FoTr1hJeWJyFIA4O+cLiSJN+2HrMQ9CW48GF5agIW4bxsaz9fII
oKMFzfrzW+YjS5jIWZMoiow6V31M4xboZm9SWUAJSll/FsXOdCyWstOWU1WxzhFYFaN0Qcn5Rokv
z1shHe/+D09cHFDd82TUsLF/3qSvCZAY0ZSHCbWF0AUg3wjZSC++tIFFPPYhR4Kk69jZADbtK4Rv
OESI0IRxyK2S+AdJ6OoMI0NB6A8r0TUUmKfFSKV5evwgCtZZorAwbYCtR5Uee7nPf28RMyoRoAYQ
Lvq2xom4HEk2fKbumhbNUxQtCcR13OK6Pni3rDNtpGIgEOMnSN3AHd+zOGndTL0H4zKr6ARfJtNU
8lP5DH1atYs/juCm6Cajl6J+SihHoTPuAXelf9W1AoTWUe4Z7Gql8fcj6dxWBvH9vVL5a/tZ9SZC
upVGniEPyxu3KVgowQPa6TKTT9ntRQBXMTfubaw69NfTVwF77LO9Cx//lJ4IHImT4O65miDp8SSS
H0eW3/cCDR/JUBpTBa67WuskIFPXvakV6fQ5Rh5uAtveu7ARI9PIu2TL4tNWs0WrDooHP/dCoOf3
cbz2ZxffedVclPco9dAzQMv93kHk2GLdOkVBXTrifLvoDKdvF15xrFM956ajW9TLzo+SHlBJaYZk
nAD3xFREkMk3ZhRYKSoNlJI/YhtZ1iDy1AwQulh6m2BVDXgn4GugjrBWyM2aqkSyhMH5mUZo397h
TLrpqE9mSXiL1vjvamn6p5jaEQ3ORs416SU8M3fFS/d2oYc5obOz+RyoILhEhA+EbaMqGw224jbp
wHN+/E6WnRSryai0EetZGagkgG5RMLKflgbEUhC4Cq307YNpYOS1cQizza34Pd/e4bGxiaYncNin
9dgDxTJG4X0gNjqKN1kEJeEVAR9ntIr4LOUkdtvwPsNSJb9XCUzeNwSBc4r94cqb+Z9ucFlO6++x
rHzFwaluVPXYAGhMKDTzmA26sWxgCEoTPCUzbmIvdxSDRSrVOybMpLQVkdCbJOi4iAspvtcNAMbC
5JN7NQCfOyzqCNU/cGDu+nuh8SqCMUQ0bdflfu35XJyGDk5Qssga/wwAkH35gEqCbh7yUt+WwDHj
+17ZFtWPc73NPfAm1WGkhQn4t0Z0yuPz7XA/4CsIyhZ3qgSatkkncgrvk5OqpaLzv/KM5368Hg7x
cScnBJXg0NtkBchVDAsRWhLaxrirexs42MUQ31yZwkLORJaogzRZxnta1s8Jv/6wtyX/QZtITc3/
CbSTHMje4qIrGprk8TgHkceXQh7sIeAHl+nTZtPPHhDSpvwQ8cI0fgQrtrHDJW/JDgn8JZNeIfm1
Rql6wz8Po4tk2kfM3xqLnYujSNfaL0cOop1rTQpWhoM3IyMGtJXkP+4aTOjeIHvDUT2zngsplPOx
50xZymVrQJfQg/WN1C3Np4G5kjcdqFKHo1ryMtGXbWBthbJJIR1SfkZ7JODBSzc7NGguWSmNnyr/
3dqCGI/nLmFzJX0hafD7BNTLJsh9tc1ybeJPj8MyxT6HWDeMC6f3aDRHfp8r0Q6AGf9TI8/2glrE
4c66bVxyaANFhh8aCkwi3Mb2Rc8/Z8IwBS6SKTiqruQMmiaezEwCZjjTQQKLDMmu3zIwI0EMudir
SL7hjen0+SiyCCXAEpSvONM6wNGJToRfTnCLEMoc8AYa6E7R5KP1RmwGNi6UOzQbS2ppIwtOdiMt
OaTGdNkmcm1ZpDkhucs74ozIleCjh8dnq9LY1jX03ZbVD5mf7VHoSv8XhAQO6t2b1/gbqFSjNg9T
MJxeJbJyEnqB6/tZUQ8mqBnX74tzNBzv/Kcxx+JRVWNNB7+egvNALiB7KydSZEGYVGEaARtWi37o
ubs46vpIJR7H/8r7J0txiBfO7QjHGmKE/7MB4wlgKAOLfvErVKcF8huWHQDcec0n508FmpvvgLfe
yuQ9D2W5E/inBDJNWynrTnGUhxQz3VPbcH9YlFUDlmlIBI5hR1US1ASyw9N2k/6GMQ9clCRn+vf/
9V+wWSDbR6OPeYEqYZTqFcGZt6D3YKD1rN84gCKLwETqt9srCjcy5rTuspqsNCclxq22l6128fWn
8sPpgZvOq9XpMCmnGIf1HMu/wa1WaXm6F9c0NCAhbYoTJX8sWosDaHb5AcLEl3RXbCpk29n8wUCC
Y4kVDO0ejiylSkeeQdLdoLUMu/UQMG3OXNsonPJ8QAHqXHUHh8ipxec6zj3xuRKAy8SaNiQliHfM
Lt3NTHu2N3nf6zQFZ3YsGruDd856izpr6jLBoQ/vImj0ew8AnIOROi3liGWzqRyu4Txs211fyUJS
4dAZM5z89fRpx/qaIqAdQzc3yGXw9zdISaTbDQGUjIV6FBPG3lYkajcZqli1HuYgQXG1GFKEU21p
BmXDRGfdWGZ3XyD/E0TI7YOn8VZIK1o+th4GRe18hYcLcdFHimRV25R+bTGccG5nRmTJ583S5Hqz
HRqYlGFg042Baez0GlGZAxCIco215zIWDVN1GlkzrrQZLPEEAXcCCMFXVgSBzSBoonudGJbAaCNd
OhnLxqRlXvLZDquts/SQnKL+DH5vzOAeCOQggO8tx7ApNkuezzzcQvxLMvXau16sFbuSjqiXvx66
BdbVFQsp+Tj6GgsynwX5mzHadGmvHRkjsctLLT3s4vR9i+2m8Wp2fkYy6YIutMYr/204vp5oTDig
ffybYGIjNL8c4tE9AMW8oo/afg/JCSjryxZWRucg+qeRr/KxEMOg+tVOh5b8c3xxy0kKd6vcUluV
gL9qGETj3FTVUgAr166cbi4330TxWTKXZxs0yIP9XtZLViOwQvIDCY2IvmIGsZNruzDFoaYNygHq
09aC0rr7Z+BnnrTzx/I92gTvKWqC+klRhGhHwSoietrwCavSRooXzFuGNYbKRboeHgadNpLq7QFG
PwftDS7yCi+dGEX5Tio0pe2ytoR4NEXQ7tkDFafY2Pqtf4U0DCoAPh17wpp3XYpoko1glbQJo0eE
GwlLXHZPRuV24lqVRAIRJcvHeP3ilqRipdY1JzGsp2Oo5lkycQ9vbn2njPV2nKY1xFn8BdeeZA7n
qoikfrcIFSwJ0ptTCDLkonB3q+40ee4Zo6VLViS/C2qTQJWvEQo6/7BqDAvg0+Jvwg0BqCtkKadF
12aPPBXhk6fqD2C+s0Lz6ZBLEjUQnG3oJfhpFziPO3Mf/a+NmvmDt5LPQqrAHYbbsNg6RLVUcneD
8VPMCKpzc1OTd/YCglleGIZZsuD0yn8787yfEkKSspOqQEHMT9ccsjARi0d1pm9JJGghPdT8H0rZ
bF+uz/MLsXSclQnfPOw/J7mwqmSceNfHdRT0yTGHkmB5SDX9gdrWSBZXfMTYq6DTgA3Sc26iCTsC
k+C2At81g9hDWceLB2h9bN5qFrQPbIo+/nITKHHQPNU+w5S7smReu2No/REpveQVI5V+CoBfsTrQ
vwlhWfO78u9xoJ8RFV8y928LPYw/iZe6U+9vWHrysYHDtDKILDlyEWuO+CmGpAujCkb2Ppp4fuAq
OefQl256uX9MZYnYHTNtsze+NbuLLbB/zNEiD5kcbpTJV0F+8Z1WGuNFlY0vt7m2kAcFCT0fUT7/
Ym+jgo8RP/NzH8FTsCnfNSdYBCxow/VPslRqhkOM4yWy2Knwh2D0l8WpuScTc7XQOMvKW3SwT+DD
IowsW/dbZXdSxAtG4oGZGm3TCVZtUKWDHAcOZdc4UKW3+ihAXqaoIpaYUmMWyEMc5a+uTYd1ABN1
acdUpgVfX0qK9PQqCc+tj9ctmj4Tc2mDLQkO5tsr/crf23+RgEdljtt9exIna6MmoyLdAcaPhPeD
38mRK0UBs0/Jj6PcjPvFSMBTBwezB4eS1pq3r8MjTT9nnOu1TBDOAIv9CKf3/159G8UxsJkjEyga
g/X5KwC+WA6M/Vsf4XfuoG++ncqzrFNS0DiCTuk/yVeJx6Xq6rzIOcf4nE3kNKGoi0658KwrJdQx
eDl4KAi9zkGRMbwtrNCMdk1Y4x1e8C/PmhPlESyXULxgqPeJBxqPoFHpCTPKm4+3dXTwxbQ4o+vd
7mQXrv5eCryJRqECr/Fn6wQGrkBZz50UEwVh1sQ+7VaDYz3R7LJSlKuEvE5sj/FTFJDTcMiT/fFN
jGmm46xBGBdxM/mktuKLyCYNdbz9oNB/zJFohj35O/qyEPsiD43VAdWg6gsEoYpCjmjuJ/MV5Rqz
jMVSRwbRk6dDcvOmSt7gfhrRvTDntH3chNl6eD+psrHRbDRurZ5igUk82eXr9jgisxHfjyN95tKN
2xviFMXRkEH1TYOgTVonmDKi/8NfyXUIVMrF+TUN/gWxVJ6Vqq3TTzyUQCNoBSGpE3W1AWrjnm9V
DbYlODlNPeD09+erbf7riqJcNMccwj0rh7uI4CkjT5c/tiEgdm8NalWhnlu6VhhYg6u1X8YOENTx
krgri3XMUhTcl/IvsH06bLdYnSmW9FNDNF7bAsHu5viGWBDpSuv96MVKR316gtL85bwGJbqBihST
KgSg0p3chno6qP785PtrmacuMb3dEeAKmp4rzib9Y90QMZF9XQLqaIrTZY8S67kPYUHbP1u3GYWV
CjeMTJKkg4CwtJ/fP8AXJJPzvUX1qMnPGqH6pFwS8/wQHuvFv1bWniY6+Waz274FsgsSKcd919cG
QvqWEcrAAHjRpHlydYnLIxSvnsVf0Se/phGnN1cwW1EsW7ijy3EWwWkT9/xnSFfsCz8jhfU7oC8J
sl5qF9curt4AXy/ntI9/XbZ2m0/fMq3w0s3ooPHj4Dd9kz8KHPsP7W4vg+e+i+lXqKyUtHjPXw5I
95JvM+oT0Cs+a4tSnHTEa+Bpz9vg6t9GtwAzUjw6qRezDtcsbXP8ElOhsTHbiGYENryTQQ1IpynV
y58WvkHX211nJ0ScRrcEnX7HuBU4uvXmaUodNY4VxzbGXLzGcWzGy6D/HrTzCQcJCih6Sqc5o+qx
kn2EwqnHtMQXmcs4pbzDaRHeiZnLMV4vcFY4vZyjEpTAu5ZA0qZ/EdU831RuYPDzlfXgLc3fQgEy
QxIRP40JJYbq5DGWfzHXSrdDOvUdIamYGqz4asEFsOcB3BnNdZ64Lk56V9RXbHzlOWe+ipkR0RH+
4ThLfHP0kWDHvRxuoZLIW6VCfwIvMv0DcYi0nWqmZIPPIZ2ulxe5msCdytvXqSzS3l/pfBOhqBOJ
pqY7OFo6eDMmoCo3bTYhSI3Tgkq3j/ZQCDzhEU8LGIznX5aE0ejrnsnKz44QL8QtiH0+vBff6RX8
l+AUHuXc//ewxZ0KV2soSbwWqZ7HiNGIVpAUe+iTYhWcFMaCU+ESIV4jIkIezaLt1rsBDr8vmrKN
tNeW5BCClVTiNI0aIbdpV0U5UCQQa0ofjilQAFIbw9TVsqncuLNF6zBz1OAGx70qGeD3TByeD/Te
AUBzMuuW9xE1Rk6qXQK5VZtxNaDlDwo27Sp6Fr+z25xll2uoZeED3LZauMQSsmxMthYkPZDoSazx
Vo/e3r9PNAmTOyD9P5q0/yiqdbE/Luj1gbcKHH4XOqbVuvATaOx4pV4zRs2poiZl7fjQmJeeLoUx
kT/CmO2ztoSP3/JRVe0ngtYT0VSNcBKWE/DX0vwFrmKE7d/C8ueGIHhmCPPaBCabcJ307FXoR+uN
ZXzHFucLvVQ1NvifESYB49L7YljrSSOyF/+miyZ9mDjxOXcNMmZNERB1FB9c5j6RZg5+VdP07q0m
RinrSgtMewhZv5MVWJc4HcRUXWpl44IH5IpG0nFoeNfvzhNTPIy+uoAqacBTouhorASjlQ4hI4DD
bvPCTB7queM5k3g6N3mIhhjfJPh8RDwuQBR1fLbFwpOdx1pPT6pBQlimwbD+8hVUt6jSr1Ewoyvq
vjBdyMvzeq2bS97qQ3OMPlT2U0T39A8pWaTSxa5lLhxLZJC8ptSC7vfGX5afD4jyNVK7ORKA0JP1
lIOQlh7LxMwdmHU1fkG9lUfXqQ+qBMQLrmsnREQX1a1W2cpJNFaNdpIm86hmZbgnbaoihqXmWCs6
QjGFNhfzn8rp3RL4dt3PKD/JUilyM56QPQlmm0XoBy4Gk0RIU5h6lX6AIDJuXoK5qF0k3hfhXfbO
cHJRArgEjoAEvEtItFj+5PRy1Lz/Uro7ZRi4leDvotdHrQShNNMEh5LsPG/d6FVMK0WXEdcr702c
XWMzD3UMZDx4jLZARORVyqrAjh6WjbnE8kbTaIofXs02xttYB2uYUlQ3XiEN/BAgHcxdYjdlx0gM
drPfeKaKJVwXVYeq1jtjYl2hKZ3Yn0EcPcwjnNfcKasYTorwKj2lL4MYYCl8/nm2dOehXae5Tj1i
3I8Z01diMTaZQn7Hyrb43Owl0OlYuRBLw6iKRBUYtHCr0ytAOAhoWXcIDiuA59Bdyv1JMAAMIz9N
zxPNMTqemswyX474/6vMAcyS4YypQ4/7FSSA5HTQrz2FBRiOWlvsWqcsenr9FtWhQ+WmQG79QgOa
ce/pL6NGG/wbDoH4g1w0bmGjBJxBx6pQB4fAEc0cWRyb9k9+HYa1YNlQPrictAXnw+7JexT6qBAX
DTNTz4bHscFBAMxfRpurGjDNKzWy6i+v6ZFjyZJPK6/4nXX9LR+Ud/syq6xvsgDzgbDMk0yeEjqw
1DAdgm2t/PFR4gfGt8moufK6JITlluZcyqaI35yilS8wIZ76rgc1gvG6f82L3PymHKvhqvAnWP5u
TS5i1rUzbhD4aaCmdwizNJLkV9emzN6sAI04L1QxDcvDb8K7aLAJee33VbIUg1Weos1vZ/ImLhTi
MKO4bXZtxF1BuzsbQ9s0ZzRVdtrZPgZCTxfRPnWI/Ttx5nzk2/iUlGnUXZof2bFg3RKotb9A7XWC
zupJsFMCwxGbeja3IEWlw5MOjacjXGaIj9BeBh3YAMz1/iuKoxloX+vmDj1+yyZrDbYNH9/Q7MTf
hiNDeF9v2yFOvpUi/MqvfdEitMbleXSdJK4xpWth1SwatxoOs+hOUgzLWrC5ndvvPE+HtRGRQEcT
7aqAYeAlYCTAus3gpkXmNySgNXFk+wqmxMPtrv5SKVcYSgeptdiYy7qvfpVha1yWgnR47RGJfOsh
QayyQUqL8rRiXtbrsGudYnELx5cKlbinl8SyVYfTWnECgN62DNZ95iZPDkc7wedU1NTIUY0A7IQ+
plLEp0hw0mbH5wRS7kuNOUfWMK5PJOOwcPX6CsKggnsmyvG3b7JuNeO7+1iXf95jfKeh/VO52Ef/
3L0R3ANGdfrAT1daD9bR/KnMNWR6KRvCdMCKYkV5BB1tUCLJ1WBTxNjlMurqvmRGK0v6cJwfjFai
tM66Ilt28zObvhx2d+coqazcfB2QvG8sBH/qvFSL5etHTyy46sxkB9v1OUZKMd0hSpR8+/QY+JWf
SuPNuhJtsWoeX3Jdzj95zzBnORD4aEgRixiiJszlAgjkCncw+KpQdQ1Fco79cQ2Tc+9KdwnlC8rt
blb2zZ/2s5mr4UVasae4i6xmcyKIIH7Lasllm4PHp3DU++XMJthwTyZ4y3mvAs4CAhzb0Vz0oZ7N
Fiz7sm7937lNm16yxN06fjCK9OlVzVMzhIy9CztpMl5H1W8vW7I517me28VyGjFJ+xeWwF6Hgv4N
kvUuH3yWP9Z4EGIGtp+/oPb9AxQf3Q6fT8k76Xpm3UA2s/MN/qkowBlAqWypkQs+8ekja5BsOPht
GVwiklO03Lz7sSUXrrecNj+SO5GQeMTySEQ78qKl+aWOoODouolNcxzN5pUq7ZzqiXDsnC+0zwsH
9YEqzXoGIAdfwAER7NT0KMcB15WOs8+MstI6oKjr3jO4ckKxmuu5Ywhu2wMEya/s/iQR9zG2JOuG
+1nf+Iu6+hinSL7sS+zLpKB7QAntHmCI8+wcpj4XvC3YMKgZiIpYPPwhfFkRvrkidQHCY5q0owvt
EcVFkiPEnQZpBgQSvePRCxXG5b8r/KuMiUfPfNQfzn4Yza5rxDQuIwCK3faQ5Lw3t68Ov6e5dSE+
hxoOXe1BazlaoCfDsGpvFmTEdpEYpHsybmxpbSCeR9kshZHKTrdzFCIkkDVfhBE79KNW30jjlU2z
23nfd1TTzvIGjYVaU9cxehK4Af5A2grNDTXfnh7q7bxQDfMb0BzMs2qfF/U5s3sECr+eIwVIcy3f
WhA1DJmNJKB5wo3dHrJ5vBucr8+Bfcv8pIgHhPqBOnRkKuXdWJf7NfWmOhgfTYqRECpzHhITJHZg
8uGPwMCOv9+C1E3HFgp6k2HPtYJUXAUnRLOFIb4IGoovHjpHVoMHak18BBfsgzWdJLUu3llRD07n
qlzrwDejGP0fH692w0Kin+T1pMA9j9mEI6PJnT6qWN3FprJ9EsqZ0WDWvVR3b5UQaW880Mqm9aT/
/tDaO9aWX3OOWUftOZswDylIHpUucKx8X8nyW/zYnKy/SBCcB0fmC20x1H735zc1iI+fshWFulgC
SZ8CR7LONEXbbsPbpeNrSACrnkhYBzBZM9h8Dcr+wX9FdtBh+dWOBgnmePpKD/1JzE0zbz8btYfU
UC3y4D+InqHiyrEc4Eutn1OOymM6GvvthRqm9fFTwRmiOSwXI/4gwXjT6s+MZiQMqHU5B1X1Fnx+
TyyAAS1YJCUWo0QNXKg5vkKEc+hyfzxhfOlx3bI2Ai54bNNBYUEH/M+1hgu5w7CcAFISKwTeO/fB
UpXd4rjaVTiIQ+J90jq8KpXpv0uqUHgOd35VDP2XW+L+FuOVl0+EbIEdY61h3I4ad4SPbrtH5gRx
DA8Yh25J2phXGD8ISvKuX0AEPnAOWk1lErNkHSCnbfjV30zzh3GXv+MNMPC5sq4sO/dbuLgut/El
R+zTtJ0u5T/lQidwqTj7iWjAz0z3d3DWuXgRITFoK0GbN5eDKX5HzJIk/2y+S4qAhErsBWDQfax8
UsVxvFmeOfRFqpMgjLBfvjpMtAEH53cZqpAjJgrqi3PchGxrCoVhaO9ZHbcAMjqmLA4RSfPLAxhv
O+te2qz/Frpn9cGS200dTEHq6nTImfEKBMtlRvMEu02OHxnRzaO3KDFL9Uir17yfrlhOf+DRQny9
lCFW07L4qQqIlqLWlcmleSqidR5+4COSNBzq764HYQoLOWNUvPwqSvWf6vUcQMFT+u2Tz9D9eIRn
f2/9Jc+KrLKYO+BvMBoo7lU3N/11yUuxoTu/g7zyB6pBL8f5r9u7OZ5QkNkENDccXbFBcy1BUHJx
mJcaazdaAqWF9X4HynBwRK1sNkVZawOaP06JGG8O0XehZHCwYnU7ORduuUQpX5iZEm4Knbppb1RL
COH0L50Kb/FoeRxy9JWoi3FlChGzrcD7pcjteDjkvJN0AVnxYvdhk0Tu6tzxX4thmxJt0fEFz2ON
wYfca7F4vWa2XF3T0MzVUgGdp1lIety/a6ciocLPSrR0RL7uD8ORgi/sU1ES7PnywuQufr2Fd5rb
qAKR2dOXVM8j6HTjQC1mG1iI4+1b1YetqnFshgXEMc5FWdOIBx84Z7NhRG0zBofXbqTTbbtmlggS
1du4xdfKDnCqUNxMkRnnH6pcVxYj/h+28uAZdpJhBH8MjWgUs7xTboZH1rMQH6VvtWcqdF4G9ECt
cl+RFpT1KmYWiMGiTiy9YRaNNNQp/BBuocMGYFdZED/G8+PgsgPne/NxluzNLdaTyfnlsFjed0vp
oEEHD7lXnazpsnUwUFxT1O4gVt94oKUlwsN9gHdAFOzIPo382rxJdrye2rl9vkVdzKHlhYGKkb/q
rw3ziX86ocUvxd2UmO2jJPi1E91Doj1jWSoFhxinvAJ3bEh7vAa0PoM3AMeYk08udjqGn18KPsb5
jTsrsaGR9CvhcVW7IbTBr/uAvirKUXouC7cLemUWDMClDmxjT9N5LbYyStzkDamVWvUdYsYOrf3t
ZkFeRi6NudXesaN2FoId9WXnVx8bPY1hOndL7TQ/Cokc3GmLCn+RZzxoXGMeEeLOJQtJg80CxBqy
G5eLmTCNo5r7ECvoIkbrVSEJnTSJ7g4acVm5nSR06quxzm1JSqgQgNDVWeTPbYbIQHBkA2EGJYdL
3kglG2VQkVvH/pmh3uMVm/gWyoAWhZbCF0tps645Osc6w1fy/vAp8tHdHY8ChIqmCCYNvuDLsWdn
rQRz5Nr35oT1yhO5aWE6awXK/abwB+Sz5ISKPrskW2R7KjdQTs996tYdNfWJ7yDjcS9ouIyx+2iv
DbV68UpxuEg5TDHZVmXCaEADsLV1+8a2XWjYxfjJFAixZQRan1nj7MtINtkOtFKv+fJaEAHqhc5w
9hJm3Y8TpyFUAhhJvb9VBrlIP8vmoJIZf402fKDxhd3DxCBQ4btMyN7Nvt7rNvJtHOJxEZWyIf7F
hcFl8vvFj51CQlgdkgrH8ivsg/fHTv8SvqlcKwd6oAOZLq9rUTHUUvKHgslrGkAEPorShEIWhitw
rbmF49ukDCKX6FMbYRrIwqwJ4xpQpAf5pNv3TpisBgwrGVWHUQY4B4phovVNrTeDfUFRLzMtFpYm
SfJOFdo4xEg0pbk8s5mw5Byjq0ryR+Q8k4n/2wH2HzKEBacYlF88huhMSAtpvmkw/A++c+GYTryv
wUYImIVeW43an0B6aL0B5AvNIKHW3JCW+NNzElRPhIiYMqwZZsroV82EqCngYX2MhWGAxkq8g288
DWZwvewUHBCdg4XoprOH1KPQ60KM+9JcmPqzhBoN9osPzD08GetUFu1A/R76ONgUOBxQQPo60ZeH
mKLam6djOO9UesSbl2uD9iwKNp7Ufz38NQrRu8SW8e0ykLp/ma1ZawAQ2qmx74h+ryXVjSSS2Cso
KUtQBlz5JXk28F7yHB6JWseZq8AOeUHpLHYZc2wQaQczv5a6Ycifm/V1Ljp41lnSUxBJHqz2gJfe
/FQPlYL9uCR7BJ02rUisJC7rpneLj8mtAwPa5RyYhSMad8xBqdGM4nPp8/pVsLoSDWmVVbgKaAds
gkJ6lvTcUfHj71cNPfJuDYhdHbBr6f+tcjaKGrLYi0uR2TMQxU23Akf6W747Yg3tQnrRYaYyOYtC
u6ASrNBJNEgBDMcbIL5dY1sveMw49NSiOffGYyMpNOawxqhW1tKSZJxvM1A3pZn9CXxg4biSNWme
XxKO2pyAc53obiJF8Jhbn/9Gaj57OqH1YhAtOAIqo8wzl9vaMMS1AjPrFElyuob8CFrNA4j38Riz
oMLL7Zt1Q4IGk3u/UX00jD3Jfq9EoO24BfuXX1/8Siq1O8TsHzF7u72mGjAsB9g727c8NYVCe2XR
4+4XV5hFqD/KZYX2z4jUW9jqI6PxEtwF/ye4kTBh+8kLSJjvR8j53PciQlbZ2daEnCaCckK+uwEx
WjJm5SX/iQWfZwVCYHDibIR6Z6rQsNZGY1hNg+gqGc6OfVxrAHLNunNXQ97G7Gv1tEA9sicppeyg
qV/ZlAbKieGHUtCLOONqRCNf3pvQycpkRVwFZFxiuk6YKZ1tSTPBvkEetGJ3ED/8kG4e2TObAbBF
qF9Q1VxfEbPrfnWLOj/kgnLp6mSDQtYVIZeCiFR9n93MZsA1w/EZqDVcJrAItuo6iU3zhyy0QstL
8AJr6IacHe4rI+q0uZ3Tuxy5zXNs2E8j/dYMlxIMxWtTeR+HK+IJG2XV5D1GH+6wR175RSdEmLeO
FR0Gn+VDHRLXsLhroR12KZ80AxhoRysPiDRBFYkC34CSP8dII/Eb25BsVJgc9mVn4l2pAzMLZkLm
P7MUtrg+ZXIGJgCpjgeGlTE0ZnzH6ZDybi45L/0AsVnkmvCL+OnaWOy6fEmb9p6rCyUGVm+YJkLS
4CROqz8/ie8+zRDTU9kAzYVCAb3n4xa2tHF7GsdzN7/ce6NAfGit4nFK+FJMN1wKMAjQHO4ashZ2
iaxL5bYPqTtzwHYEQ8vJhwn6SrOFIKUqzgdHuD73NHBwMcWYT1bHxjKxvGQBEd4Q0XNDgV7ZEa1A
RPoa6SN3fkEx47WG0/Gg8yo7PF53jBFk8aeHU4xSh4hat+cVbHvgvdAUVKXlTKWuHZvtQYsAVOlO
iXxR+X6+znrxPkBQRM3NVXTg/b6wjU+e2aRCFdRreT/yLhT0kDibhDI1l4HkNZTSjs1hGxoYmC3c
e/eb0r0UJf8yq9GQdrOuD0CYMMnPw3nqvojrFrKujox+/eDKtX3Sy1Q+z6+LQHXK9UqnU1RRpR3Q
xKOhPb8u1DZDFPi8Me5hZ1CxNQapy4v4b1GnW15AFTooNI97Sow1JMRaAcfDgWvWSfUZUy8l91WX
pNd3g7/CbcMK2qwe1wA6OnwQjJpqz/9qLU69XFUuyBiMJ0Hq4XJ/UUfvpWKodm4fElnT84ca3deQ
S46PZAoRv2/2GuzYLHw6G3kEURnIY9oTrm+nba9QcOT8PnFECG8PxrotwUeHsO9zD7laajazDqpO
HMOFxzPDNEuS11xPsW8Qvzz1FH0vBtl58Gx3BFf+0Ik2cbDfWN9PdiTnA10sVuRZA1M4jNLDsdDF
f3E7O8XC94CEeIIVcuj6DCkTGDycTCrCjiduE9qL/TA9234zwjWS8/71askkMy0VvG1FC5M0ElSw
aNN2iQj3TABSfUbOjJS7en/6WKUPjJd4CRDw/9DbfxhxJZrfw2rW2rKtgNKILHr18lbZ1Eo/rHTg
zcvufg3oAyi4wdqFi2GO5eSYmo31AvfmF0RSHns6G45zOaE1OxcH0b57jcBQu2drfRkiSOiDzN8/
+waRQa8VgqBpQ/QHsl1DP8BAXzeVx1NiMvSlV0p7aQQT9CwdXiJffsjePAD1IaCRaa0UCMQzsOVs
0SnQvnhYqtkz7XR+8Bfl0IpyU1oSekbySdklKX8AiwXg1oznvdXYIyQzWZ4k68gZBVN/cggF7MeZ
ALNLKE+iAiZi39maIGsn53AeAyqZnqIYI9pRArZDYcO0Y8V98YbT7XTCPQKzG1adBlVUERXlB/4M
n274Hsq8vOqlJTcIHAJgm0Nc+pD9xfHxJLAb1u7MXgqvhkflnKQ356/ic38L6ol4Z5ShuIGMRlnq
JfM3SqGE9cJxXKP0bo4KG1KmVnDEv23ETmUGECpVDtXdn7/J/E6vOFZp46o08NNJ4z4UxhN6yWVP
u7FCzhPCPC6dOPjfH0bnGvGvHG9RVrUTHd2VvassnlwMWWIcM2mMznaELaVyo4srD5/gTxFuJfbY
xxlluKkjTdQ4cmIARRwuOdjL6oangQReTbHXlN0Wjq75IQqwG9L61VlBVR0ha9BG0AjDmoEDt228
2IB57DRnuDcW/NTVtdNKQW315ckuOwN72fM8LnsA7UHewT688ZMQAt34h0gvQkf+pcHxxduBuEcK
jaRgx8oyx5lNEq/xaJzWW2mlqyIYEk0c1EfJu2wxo7y/XmXYPOgDVCOMBs1rNoXmLx8nBu9iQ45I
0M7DQpmZGDitt7Haz6T/wqbPtaV9QioWCu1LQxe6zv6L1IcC3zPLsVdmeNneuVIfPC40/x9jG7x5
9YNu8QPOsfEPZlv3S54NUoopuYZqPTkF/ojAdlaF9CLrS2sloVqloVXWDUpB2ZBy4P+ptXXtD9KR
brt4ZbV26w5dpMrsXLY7qafYVdhEQVjS1HXYSYjnGWzrMdGYWFEdk9tXrGdZ7sOFDMxcfdZPP+OZ
Zjd8EdPDEztkeFVQ3OlfT7QwJ09f1kDjXo7D4M/B9pKlDX7AVp612MqQwqDwqrI7wJ6YH7TBEKSG
eOz5yK5B+phK+udShgfjicElh0Z7cJ86H+SzLX33fvgMpTjsHIMOx+jyplfj4fIC0y+zMec1Hf9s
8d3FOgkShp0zQBfzti8+snUKlrwo75ng6shusqG45HGxTJTZ5zdfVBeqpSwrjhdhy3jjr7LxfOb1
YqT3Yy+3hoFV1puJepmubYByR10SnS8/XEQaCvZxa+nQDTkNYTMuaExU5rBSKGMextZdssOr0ZZv
fr3bWLiluhW7f5GSKGWqNpfFGG3VCbO4KBdHNWeIFLkLcQvcaIrGGNUMD5cgic69pX2pWeY+RwlU
WtTDMBCgnmvw8flR6k2o/u0HHZyVNdf8TzMt81gh/mSxgXclgZPp9cx8MvNf6uZrs4or2O710L0O
kj9nbpVQa1X9ASjGJmM5b7x9l2o+0beoiPExPDYNvjwk0VFlM5TMVinptzTjYBeTDOgm1zAhwLft
OzovwI2l9oMSM3gmC/ED1K8+nwE3s6Ozv1VXv6lJfahaXBCK2VPqU5KGk/XckCWI28lP7NsLGiFW
mco+aLMh60Dw9EakF/z2dsk+b9rc+c896NTTNEZA7n3b1/LQs9c/ARDOkxbG2M6HHeiiTccDn6Rt
Y8u1JbeHvehAIU8oXHlnP7kmJYxFcRPwy3pUdtCDRtQ7tIqNi6pRCt3dJg/FOKx1jOXFnf76PrHv
QAd9dzdexh+L8Nmuyw0scmx3HB9aPgqwhdw2VB5Mda9owQim3lKvjUvfwMftRe4Bps9TNcFzAcdt
xZDNXKqCFDKJXKxGt2mOvOgb7QliOO+dsKQWikA3S/lz3mY9+pPxZhScpLev+cWo2tBaljw2S3sL
61CPCdLjazGOJ7v8N6rP2Os/ayy/i8bF+ex3Yh0FyDKTQY5quzfYt+G+XZFuE5rwTcM6XoO+/Duk
UzRc5fqd7cgQXDqIsuvwqDtMFK9pjwOm1/ErbOMKQdVXo/t3wszqZV2nZt1SR4f3JMDGXER5VIY/
rkexRjYA5V910WT29iaU1QjMg40JvKsegxXbi4vMCMLBvvsXone0tTVgOJ+rke5R0wfe9Ap8bmQO
MuLf66WOb71+QPl7azbsn/l6fGpOg65RM/xzV73sp4yGKsR88lk3mTIxGt/jMU8XcrS5myKQliJp
mLoTqtTvPixjVQpcUSydUKH4WiWODC4Nb27lYkK807yz2SNXV4iKO4XsERg/c0YV4lDG6tmnt7v3
UBu7fRNdwnP19PMehKTFx22XDov2iTadWDRwk1upaL31ohVILZtMTnekp+TZ15HeRWIn13YVYwOE
NMr2EaMKRNFrmBT9NX0wNg0jYbwOy/lzcQMEMcq2xtuHIvulmsZBLFBGeA1ClVUpvBd2zvYgIezD
ms8eZgD8nDzWZL1Kh5R0FrJ4af+siFOTPBY2vTEdVju1uUPrlU82cII56y6pDvscUSuNHs/GodXa
Tx9ErlaYMcfqM6iiwAohwnPAUiLImQOkjYPocjOpJ0qcTgCviVgb0HyTdADXGEzInRQ/tL659fUJ
844wuDM1NBCVI/UFKqw73dby2CcMD57IuRlxFy+26ZHKcX44PlvVZrdcppNg4tQil9UJx8yoXWwp
YRQXSABOx9twjfPP0fGHqOZ7zdFR5nYm4QFQGMdLGpDLekofTodsD+P2Rt1ZQSZtMWS50a7zZl0z
LJDlbKUB5dshGmcamhbnc6plkgF3nf+1uOpEpo3F241aF9SGC2dJCIcWyeY9EubRrPIUQ6zlYbF2
sXAiSR15BXawz0V84YvD3F3yi1P4Cwe8xDWeemGl0fFsv5wd9WWoo5AmSygXk0zAdpR6u9CjWa9E
bss+JzI9ULh41seksGR1VTNo3jIhmnI2gFhmKchrdXsZ6J2zrcltQZ13YGUB2pxoVGg1QRBdzrOs
IBti9lCihayjAWcVZ8ZN1ge4+nQW6e0KbDUjRYxt//i/Wc4oZM+HA/LPiRCeF7QOzXVh++Ww0S61
17fTQN/jlJrS6QvFaftVN7CVIzc0twCHUKjT8L+d+icwfOdu5xczrTO+YBk+sCQvrwHkJ2pzfiy1
Aoxg0KHL05uBzBc6PPtps2atw9toGbM+8W0cQVsocp5A88vtlwdYLh+Q53pz7Go5jGIPA64OmRiH
htz9y+dKZhjJlT486IGvcFQe+6r5Wcib3cb7tC75wZrMiZTE4mkgeuVN/I5t4L3gEiTHIaH9BQbV
35uBSCCjXxw7Ner1DwGuJjafZwiuBIP8e/O4TI+cGFR/QuMK/ZTfOoxZn529AC7JnFRF+t08921f
2rz5BfIO1FBS0iUR/qbWKsF5yG5888APErcobf9hhuOCyAfpzimK2CJseG8Nn2GzSYATi/uiAm34
aLDnqubbJFpNGGRT977lALoM7lA3Gpj/NLxExo/4eRTh5vi+357GSirxFBBZLckj85kmAANfTi2c
GkW/NnOsdOW4LiUCT4TL6zemv4260w/1CYH7dpU6Mwb6ikf4vy8vvUBzZDXDI8alacex+J5Ql39V
aNRl/YP/VTQWw4vwvUpNS+ufjTArBNLc1z0/l0zUGMyiXhwbuJnUFwC83qs0ioBkUZUAyaF5xp1p
j3cdWrYW6CEtluFjQ35QPzHmZ0NhCz9VG8S4UomyfbTO6BFsX0YC+hMnTIW/TPERcl+Xn/va3kI5
cA0K0PMqi39H2Ik4I0PREBxK8C3BCeiY5HI617R4T5ZuJ6IFqkT+x9lbbwuNVYH/aBhlZR/kp9g4
KEcAR29qf2FPtwr+wNt9YGdnp1Au+BUiTcDpusvKHSQaVm86s1mn36xZW9miaXW0KitnMx/6jyha
OuvoJabdXbvVlsps6Te8/5/54mwrjiwyCB6uwCriOHL9mk4MKxuW/y+XjcyNELypiCS+abi85B/a
N4UaKu4RgGSqF88TAmju41Bu99NjET/iAaZq0b4lwaGjw6VUzb1a94942bwnJSFLHBmxeel/LFpX
uK/+fSbpcj0uTNS+Rifhh9jW6Haq4hAQg7lXEcGqQomOZudxsK0JukWYYRCeZ8E0EZXEeiE6wyYr
FcXNZyaDtQDOzwD6V9RLNnvqLl3Ud9S1KU39nmvhrefcQixSfYvCfTct7vfM2thxaytfsP8hWK76
0XJFqGbX0w6YwZjfXrxzjNQykVMbWMam/TQMc7UkGaRxB2bwVI0+vxaPSSfQlpysHVCfr7p45W7m
0/dKvnNpVJPogg5Xml69eELlhKMnKEfRMQr0fHbBMHM7lXFaNukxI0h1nPcvet+OeVSpBqESomlV
w41a5VVlWBlrkb+CSkrqzmLyYxUEMKnape+1e6QGnL0OX3uQ9AJdt/OPHvapyL6Pd2KeYa+6wcYg
6v0H0vtkrOpf8tBZk/FKlcilJI3Xlkm7VO6fejXSkAQU/c7Lg05oe8ET2yiJ56+gZ6XtBCtt0qdn
N5u2fK9rrqF6ybcsXB3fGhAVdGnseg5A280nvjULbS0zJQ8HgGX3G+yiQhiQ0mTvWE/5AyKvIsUd
2B6HvkH8LntL3zbTg/kmcsWBPmY1NbutXQGCj2oRHrcitF06s2Fnh9zPQIIyDYcebBNKN+kNIXVQ
Rl1aFuwPgnF6f1veu/lwRTNCLr9qmjlFpZLDI9UZfVFXHpV5XfvmGlRh+2EnkXl2/dVwnUN3vXNI
eIeH0ChO5l8vqCQgXGTd1i9OWPuKw2G4HsIiPiNW836UDHv7/aRwz2d2LKmRzRUssFrlaQKTX8Vf
tfcWxoL4fDPyipODPeyK0n2m9nW2Y4/woov3xIcz3ZZ5dP+YOIYEeW+B+GmR+v9UlaedGqQRCnQc
S1NFasckfH9wW0esFSfUhV02X2Rc3HD7poVnm+5OoahmHyAqf8ELgZ7ZPw0Ie93Kd/2aTTTiT7S8
vjkLU7bcudIk2deFMXFLM9eOpN3joQ65BOwhn4K2XsNdtOUFoK+R+HOS4neV8ikJewfsxOH44o4b
pg2Ny+84PIcv0oGzlXL7+KkAD9wwRD9h3yDSN/w/HE+k2uk4HdiGOcd6WG1WCowA9tVwPiiZ9gqf
rU2nPzXGJ4akfBAsia0No+V0cY+zTjBO0Dpgtx5Wo2OnptRzcEUJw6+pOrYN6E9Ef1xTiTvP7Gjo
l/mPE3xejw6UZkcHYOwz19SZAgagDpdLBPBj75trgodx/r7SwrQ7yTU6WIxLhSc9b5cpiu6UFhp5
/GTf1WGGNLb9OjHad7qUxL85dr5GR665SkCfB30A3naKM3xXQrNBWdnbqBqsSFfRgT1cFCJWfGEl
icX5kop/ac1IEN1gQgstUMcTRmjJeetg5abyMJNCxy9eDKiqIlHoLdvUWMNuX7N/up+Db3NDWRaf
86mxlHJaWHRRGVcbkt16OK2L1ZdgjcYJV6zmez6TcmvUN5Ynp7Ghj0pHKjFvgiCyxpnP8IOxU+qS
8qXRMcPAX0y+b+HSDMgiM8Pbn7dndaJYZD1fNxIYBenVrFlNZAacDBIoqLDbS6iYE8KxHjS7QmkA
7vVvWYlSYhzP3BLi3SCYeXUfyo7wUjLCE1EWGDjH4BVgH6TJar1oaS2qkMt8oW/OyFBTSqQ85amu
o8i1g294UUE19DZ0K6Kzic9MlaOIdB75GFYd3FpGJPaZAdQwLeNbtRCAcnUZAyA4LYwN4As4b/js
0znDUbb+YWMKKWcH2ivBQmSCNRj+hh1c/i68zgvbyg8C7D8aJNPXo2qsB3RN/vDp7gnQZUb7ABG5
6G29Te306hd4/lVd/oK70NKfcgnWTEiCOUr4MnGQsp9/riOeMKrvhi+bgqlWLHkwia1iKF7MYY+Z
Ze2oAy7c5Ufo8f0FlmRrORsa6+HSQLgJRVsk4YfvicutoUReHlMC/XC2+R9io/T6ngP8taoHCCYl
huNc+WJaMtTQCl3PtJPHKYR8IayaFDBpDAbVt2wSnLA9n9rYFY8JP0KfYmsJmAw=
`protect end_protected
