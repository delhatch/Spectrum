��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J>E��
�L\�īi��౉�� ��6�կW<bQAE�s����3*�]����d-/)]�������d0sb�M
 ��:/�J~�y��g�Z�C_�c���ƻ��)��juR<O�������=��V7�h�F� J���H6xOI�c�m#��JhZ�C���S��νR�}�����8��/����|ʅ0N���FQ��v��[�jyH���S�_ D�.x�u#O�{�md�q��ENk�a��v�`DU����74KR�&����RΠ�p���z�|�+3���P��0U܆
3Z\g�"f<C��1.E�a.ú���Q������}i\F�j�:�?��!�M�WJ���Ʒ�2Ҧǲ�����'G۾{~|t��?�����0U?�S������{V�~�5����c	i���r0F%W´F�����ij�c�T�|�8*�Ȩ���Fy�T���� ���Z党	 �D�KU$���e��W��O�tO+^ `:�'��t-����n�J�e�JZF���n�����e�GZ�#9�g���f�a�P���c����dME�m���1��=^�u՜�?)���fy��BSH)����2�[�8��XB{e&`\n���=�TI�R��uN����=�%ubK7�F��aL,��f��j��t����a�w���x�o��@I�����Ӛ%�=�#}2vԦ(�j����A�b�����5�(���g���y�t�QS�L����g@ﷰ�a^?�=7�s2�RU��ETAZl߁��xH�����3%���<�};�Z:�#�@��6$ܱ8�Bg~b�AY��sŜ�Y����bDU���8@�	�}ydv�n��2ߖ�\ۇ�w�5�Ĝ�wv�uH��Ek�	��\�'��l/?����+���3A2�\��.��cf)��Ӕ�$��O6-^�l�EVt *�l�=�W��`��ϫ�*���#��B����� �,���~�����������<}|�2�9�a��-O��;���Lr�QM��e�Tz������{&kf��-�֔5Ž�����g�R�cc (�M��(��BӘ�d�w�G��ș7���4n@�AG� @�R�3|��X�ܜw��\��]�z�܍�N��C �km	�u-B�@d�����I��iq�?%=�@��&IC����h�[���؋?.rl�^�/Ry�LtKED���zL�� ����<����P�������$�x��E�M��-����Jِ���ZB4� �|����_k+�v9Kkؿ�z'?!�*La3�B/��\��<*9z��U�ђJ��s�'�Oi&ߞ��J}郡3���/�ݭp*+�(�48�o�&^�%r����U�(W����LꝹ��V!w�c��E��k���̙�h�ėoR� ���`�oW��[�U�\��%�
0t�i���c 6ߦ�V	97Յ�:�8�鞢��!�2�t�α벌~X�,��B_8ǹ�>��/2��������=������^�[��'	
+��� ����h)�utc�ʇ>K����o&r�ě���y6F�ɿm����.��DPr8x���&X0I-�/ȟ��i��Z��Ϛ��qXh|� �W��h��W����6�d�Ѝo`IxKPw����j�
����ѡ�.�^L-S���c��|��cPJ{0�]��&Kyh�<�	���m���H�T�%Tt=�]�1�<�:�D����/����?Y��6�ҽ�l����Ҏa_6~,2���F��Ǯρǚ�6�����y��{�^�*?(�)���g�����	҇Ӽ��F-f/�>�SW,>�n���(E����l���5&�Gr�!Ω9��<�Ĳ���T[���>�>.	63�Q|�6�{��y�l�Ū�|.���˭��a�D��"��cFA�k,z
��K��I�`\��aq2s�"ڗʰF���&�zؐ���N?̉�u��m��y}TeJ	g�yk������4�+5��r�s���hY/~Kr�[���$� �Ղ�ؒ�)%Q/�yZ��A9��jLm��݄|V�[b�1�mܪbF��f2�U�i���_���V|'W�8G��P�`;��*�/k�\<�\M�P��U�