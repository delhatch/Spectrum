-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CV02hic4YxVreiA9Ce5+mT0Y7uvIUe/eiI67tP7EsEc8sDbykf7v7rapNzqmmavKTTd0VqYaVr8n
cSDgkUi7Zsgia19dRSCvwZ+hDx6ZWL1qPbbdA5mbLD9hsFszQ/LQetmCDmKh5ZkcH1jhKXQbO6/L
eN61diJn3GiSo3fM0d03pHGK9sPV9Q0fAs195PKplTpfONmE6+RN9ySESHX56ActDgjvhCv6uUJl
psRo9TywiEQi7Z2zdSY3mOeFhCTL3Y5y0i/E9UjZdWgZRnFHx87rbrtfrkHmcEXXoCo4NJRC8UvG
NwS2XTq7Xf0op1Z6sRDlZP3GroBmVVRDndl57g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
MHbVZGjstUTdhF25+oDS3jA8ZlXWP0abjOedudGPGL8K9eEw9bpPmoAImy7HqHN67UybFq2Lvj3x
TEA5cLkDy4u/xW17O0Qx6hGyuPu+B+ZjJ41kRLAc9tF5Z6mytOfWjksRe0yksNmOBnUgytksGZBU
IOSf2YwdD9En882Q9A0AbGfiDhUK/xPOaG+u/sO7RYf8WCClphLNkp5oDS+7Q5Wf6LJu6mvRnNQQ
Fy/2VUOCmUgWR7ek7qKeoIDAmod93666NxzO8CZWtp5ctb4WzOZfVkpuWx5UGxyWSibYJOyogr+u
nG+VY6CHr83RED0NS6dsYp2EIMS1ickxsNYSIYBiPd4ZjsMAEThM7m6uT7j6Qe9SqmrOoG8mYidw
3NpZzy2MMXmuHe+HV3grSp/G1jYPH45lJFWlS9fJyN/Xzqc2s3XDHWg1Bf7Wu49zPrTsBOm78F5Z
Q76LiP71jGCPjaY7WtsujXzFkz27TQl8R15SEWEoptExtccKzCx3LNAQj9utkO8+cWmp/obKgwsJ
WVnJEiomLFZ5/6Z7800lgrVpvtLUTjWk3GHDUnoU3o7KhfdJnndmuoTBYQfghUx1zazYUe6dmx47
h8YZul1x2yWEJPr2h/oL099xPYqMvbzOHZHJk90DY2yiLfdinBymGGSYA5lBA4NY2ucI+LulwwlK
4W92csElun+CYVskd1s7/8pn/jigvsNsDwD7Us3QD79uP1Z6WJ1pD3hmzWsZ+dXt4nKaqIHI8ppK
GCWLuY7pxvwT/pcXOAVZDhWqweYX8JYqBktJyEYV157nJAUaTgL8tdCEWODZ0kz2DvNoqDclSaBS
YIHIKlIzAFVja5G+kE/V8HBSUo8VIBqCeHKN/fhQRdzSjsayEubQ6YOQJSUW2z4srsSR3DruIzmB
jctKSRrMCyHhtliULSdd3lUAYMmz+wynJFmJbGiY/jZsD97rBelwCd00b9B8WNKVgv5pioWSAKat
k3UEcOXr5klCcEW9UBcB36+/zpFTSdbXqwPzG6T2sXwrxy632HGVSHKSgalGB8F7VBmivVFk2AWM
MV1M5waOYxM863vHFqaTLCEqFVbGLzCOzImKktZKWV66wD6R8OTmN3IMWjKJooKRsn+aU62SC6vY
dSrkkjJep4JT7ZeTs5U4Ie0aNq9pVq4upbDD6Wi7vwAAxBIfSmUmGnw1ou2XGe6I3SYJDkTWwxM1
+oNjF9gIWBVVu9biSz63nSvOMtwtipwE9Fagv1zFuSy4ozs+Ey51+ihZ9yPSaFikbHNPdsXFREwz
5k3NFXTb3rTf4QuvEaqLpMcXC7yANpDau1JOOu1M/3MQtmE+oDBlmMVmQqk5FFvRGnVl8QyxVY8e
dOb9xF3f3ocjhTeMDf8ymPLeFhycyYOAc1PgaHaUW/SiqdzfXbzZFD2m7j09mhPV3G03h7NStd5U
aYb+AcBhie801AAJjeYcr+gIsSMOYhmyDICU9XB5PK5tpfqGIQMv/ofUFFxJFfYkCyk63vN5WBid
eV0ZmBi+S1eRZINGCidNO++O/Pci00bvdk6nQh+/Kl8zJ5JQUOMKIiKLNYa8daDP6p6jQciu+y5C
dJZ7H/zRV8DSKycUfldctRyTNRf6fhRglQ1XGdh7CbUS9/SFV3DzD5bk0BU0vN3ya3hD/DqCHY7u
aVcIss4XGRCBAblO7ZUmen6k7T6Wo3ArK7dPZGNaUnpF4xzl9le0JPXr3jX9yNdz8yxCiazsGBeS
2vMpE9qX/gTFeogURXYDD/J1Ql9TCCDxcf+x0u6YBLEJDGn1exWDRTzfylp8stzYb4bSCQ1jRU//
h88oBYvOlH0unJD0ymvxgp0/pswMsSNmgitDXtCZLqBf7d+BRwwYoLX49uI7dp87FniS4LCRctJZ
rxA/plxN+9RhUEMDpPAaMdy8Yvqv4GlSH9ZjrQnteofHjQEk9N9IR6AwpiGG1lbHbwiEaBGf9qFi
42nxPQgbF1yOxFickO77YQSFH/TteX0nglfMEpvp3Ih/QNvDYqmHn9EixKnV3CHZX0+Y9aL2ObzH
9Hmw4QUvDJpAJ5YFskrpNwT1kApn652563EZ9cOBeYfMPYlUV1f8WUbhFlwFCDHEsO6DW+cRCmFW
+cVg73tAyzAd/ot/BMSTqdLIp31Ojpw8D0bZA5EAEIW35CP+peNaWsEzZks3ZQALdnEKbX58yYib
PyajiBUaIaR1EsqrTIKecUTk6aHIMBHqFh9W4r7OBVpsxMWkyly5uSb9tNgBznkwGgVOGbft8yFc
xi9a35GrSLKj7/w0pA2RZpZpB4bE3dXpGE+wPWnB0FsA67i4z58IcO7O13QmpIk8J9t+EXV2zILh
gfhD2JKQwDLtPEftM84VwddAW+1zyyYmbA8MAg/6ZQ5vykmIB/78IxFHRaOpzZ37IL+sZuY15a47
CEmkoO5nW/o20YQiz21TWvzTadKbSJFAAF7C/cwH4csew0dOivzO+dsV/+cilTP0ezwpbmCrKIRm
R5ebh1LIxHzKTBJJG8eSkEEgtBU3KwYqno2uy6l4OVL17FTjzcZGfVaqRYhq0pcCQwNM9s7GpblF
/55x/fecZPxcERJnQ+CRDI8r1gJmKsnpKlDo1ao7+SjyDmaWzihIN+6uo7UuwLs1PWP1SAufxHB8
FkuNg6T8f4Pce+zxEKVXw2DwgPekgF2ge39Esa12hcEXBxpwiPG1keVwnzSFhnYsIq2taxDZmdRB
k6WvWNKgqRLiTTezDWWQxZ/tVjhZtvks5GyPS1/TK6ff14/CvpUC+Z2hXo3DatnwopUUrWO8YMCm
1cs19+dWnTzVldGF3fqPy/haS9hH572THI4ag+oiCzyb+lUGYKlK433Jb/rAVlWaU5ExWCUlVRKk
DBQSUNP1UXmVcqs+uW+IPtXhJ/ezEwy3ETzyHXczO7YG2HaJettSkv6EVexR9eXal0gSm83eRG+U
ond4TBp5tMnf5Twc3+1oApuKBW6Lps8G4ENuVoPUEpSLMigZZ8DACLJtzxLz7Lrn4avsjkwsz70M
dUAWazhlw9T93m+8SBZ3eU90zF6H2G/QsjaL4AKNzePoTZbcRAwnXHG9y8qhKhVNBAZXErHym6Ba
jTuqw4McLo9xIr8qS7p5Xv3qgG4ShjsOp63dFijmSprIocZx6iZ+rO2uPzf5Wjtii3Q/wTXuPIDh
L9a8sWWZzCNyAkQrs+CmUTbw7miESATRm8C3I5ScOOemZw7b3FFh004t5N2KEqStPDuN0yGfhbB8
4VCWK47+jqznvh0njwqQ/pDYlFtxbQZU49JyP5/b8BaWAVudJGveLVz1ppeg67eWu8DON4qMZOgz
IAUzEnkD+bFy4wjFHJAXpl9j9Y2irCYMd0L53pdoXz0HdDl6YPPxPE7DZB3+i2EeQxHOuAcY5Y4n
xRcFHWu1mgbzOvpS6HbonlWmlg4AG7qbSQ6RAHF0pvTeDf1LFkIM2nCtz8FoHZI6t73P0qopHryy
hA7BrFmTzwMTUSiKXT4mBBeT2Q6HFo63LGyefGquNmQqSJnjFyZNmIE6F2DtDAWcHZjEm0BgtcLI
Ny0ke/bxglp6vh5p5HhBK+Q56YN1dhoM2ccZsGwmKk/26KZvUYWPexPM/rZ//rVO9IIRwFAIQ9CG
FGO8b2DcSCFyyYNtvZ9kEVgPxKvDvXW9tZ4pseFygSrfX/wDny0TrJc4KjJM5sHL2XguklKXt6um
LJ8AB/Z85lrZOp2QbTOKUnttDFXrAVxyq+sR39Vnln3i811ukA11f4q73l0CooMIhwelV+Z9EpTN
GziLjEXngWIEK25ytIOqKyU62tuRhw3+mpfKj03J9rgBea2aY+en9kkaSBsx8hEvnVbDxH4cWHgQ
Mi+c09nFIAiZfUu5zB48jEKq3yuvjC5bb4mtjySU7Sd33NXYBbkEW8oORKcRk+JWkinSwqeOSEL0
yoVPgYb9e36rZ9hb+VJ0dUMRCIoFJfFgqZChpn18olqTOom1PYLDZfFgnEpLA3tzgoRfTDQBW4AM
xbTB2felm+ylU1g7Xlanw3CAu6kCzxcKse81gWtR43ZrNy0ag7weMxVXApOWWRfcBMaAKlwEOkpF
4cPNsvLNkjxvuZq9EbkAQ/uKzxVNXIkugeWbvlExRBZ9Q223iKLcUghMh1Din/cSyB4rT/BDeyyW
AEcc34Wuq3MkGRl87/8mgaVqHwQudlfvjMMXUq0HWDQOy8t5VYf5FOFuzUxQm4iIrPNKABr7yCBb
HSeSaltj99sjNhqtKE0dgyXjyreSGouUQjru4yre+IfL/SNVJp2Czwe2eb37iCh2VCe3cBt5zhUP
fAuv4wMUWJVTS5waF0L8BiZU5H9wNfU4SoewuAs3L41LBZqoZSWT7pvPoiMMFPVSzBKmFc8/bGUO
YPtSueEGT3Z2aesvYabW3MTUjZ6tIrXdrioUBl99HPVp8Mf22I8nke0zQDL5NYEvs28Tbb1L1NP1
JqNpXOoGU7jCQCNDl8Pe1iV2F2ysYKu0z6YqK7YOTe5M6vFujqS52l7rPDWDQBfIsdiXso8FbM6W
E/KjVrG7HmpG2cLopksKj0puZ/enGHibjJdgdmhy5LQGPQHTJIQ9CKN7MzzDsHGnapuEGZrTWpiC
Mf2zcvu67ckorX8sOaNxfKHbtqB8W8EQ7hkUH+NUNNOSedUR7xpP7d8hhNe4JlJ8U8vOBruKX66k
q76Hz0SNixiuqDyl9tspbzQqZHeptLeis8BWKsWSeMeGxjE7iM94wd2aNRtFur8ZA+v73gnfVL53
OFKwKYh8An52FINNhEem5PQz/CL2DHM0Aavzr0f3ZzRU8kzHMEDRWGq53eKxp2R+RoP4tmv7JXIe
SUSAoDo/nm8A3gIe+Xd698lADV5K0nqLLau+X1NAhQkGYCW8AMuh6FgkcpcM1ij3+nKVVaLGRh2E
eU9lcXUXeoE/hzrdt3tkMmvb6xT62EsI6aY/7E4dCDPjherGqVGNHrPqDrsHIn2rhhK8KLbuyzE6
Tf/pv29WC1MvCbx5CoKxdIUOW9XnVmcRAemdveq2OaBk3Z1SdYmEO32m/FZq0vo7FH4GivaEPJwW
hVu/BUe58xFZkxcj/2XoydtOu5NClvxopEY0fMth7lZbggvobUR9I24TO3BJluCYDfuuDtTEuDgu
K07EB6nbqx2uwCCgSfRIUI9lUV4ET0oHsCnnceob4fB422P7eknEBFO+iCN2d+HgOsSp9VTq2Bxr
nFyoekugnHydN9s5x4W3XW/Sf3ZrOTRXbNCPBE3S+ZoDWCgroTNv93wg3fsv/YB4OjPT2o60j7aV
c/VgeIvPIdmBoDGJfmvEQhcGwagvH5vSj3TkIHB5yrTEH4ZJaNf9wCCigFn4zqeTgg36Ff1SIcQL
ZZd6tnQH1OWhJzCkMDEertdbCPzZpDkpvzdEp7jcsSx0PiBtvt9bCM0/XWX7ReKU2ZPjNdWZCi1t
2lWRtxfdfQnPq88eKWtUeouoI7CK3AQhL88RUY9pB6h1oLLhuCIenu1YaQ+kZWGmcrHQFsG4gD8a
riYdGoSYZWz4+dmypkNz16WbgWLRagqKVHgEcQ/yhgduWBLa18i9U1fQcZCxALS1H7xNH7op/IjV
jQdc9EH+7BToCo1TmBzBJvZ+Sw7Cz5tLOsqLlFY5aU2JET8A15qKbCBQKIpzukZsI8hmvbPXC0Kr
0YaNs4yShRQS3Rqv4ZEa6mYz3a3Vo2jBERGMdWe1P1g838lhQ1czhZUtaX8Bk4e5yzZf8TyPqhG6
3t4TCtKi+5pk35ailSdIrQLZ/bg3pqXpqZS8jopeVeY3xlIbIzNkDv6lPFJ0MztG/pJR0Y09dObX
Hnsd1KFKk7numw5rZYYd7H/dpwabEpxl6LK0h2gN+tSmqGWEYisSTSOGur0y6eCHtT9UoaceiEtE
yeC0Zs+T7z+VUVl8OxJ4PQxgVxuMkev9JrIsonZbRC9f8DVryIYptJgJFSMaE7JA5W6IUsvf0338
lMWSlqHZqMuTFnjZyhGdAYaw8TDhk+qQMQ==
`protect end_protected
