-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I7p3oV31CcdS0+JZpK7cmxyqsYYZgQCHS1qd4CMoHzeCOkUSgVs0JRBAsetNvGnbgMtOdbtPzB7y
YBqPzvcXIyx2239trWIUGBMI6KTYskWq/jjNZibImoVfTrZMhPnscbx0Hs0lJEfU37wcXVMYgS0y
7BihqHPrrlFSqC7bE+3tI2EDoHwgQLP5R4PJBHdQ58lkbZFmUyFYu8kkZZerCmtVMuLvl3pF7gyD
LQhzEkyicw+eoXTZl+zjmxTjix/iI4YK3D2zIHyk/iytBuNiHmt5EkEBoH060hRDLf0iSmQ+Ftxn
pf23hq+c1u5kcKcLa7heBNOyyXm/5J2B4deTqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
WOFiwZT5q+MJFQUbyreeLyKDF86WCBScOyHNao3yAFx5EoTQg0DN9xqx9aOSSWCuFZSRvDSd4d1Z
jXHVQ+nB4nWvtWWmwFr5BnrmUMjxxmJy5O6dksRizSCUpCnxyABW0n67JJ1k/qUkudKeJvdo2XEF
H7/yaSq4/NIPXtPUb8+rv1gcUWTPuptMaen6RVLha32Pf/0Ar7cqvMM3QDCjdHhE6NDqWG0Ra8kl
me9TKXESDXytoDqkVbj4pK+2fWYAux1pTtGYCusZaKAaqTMG8YunjigzbaaMicpEcEu+T2oLjSuS
SeeLBdpzEb2Nw0bJmQqNWuPceb60Bpl7OPMOH3MRRJ7zIAAOmoWGa6+d3oulTJfs0cn9jSdVSImM
fHXObW7mqp/GpijCSv1aa5JiQitEy/Carq9spDHp/QY6i/CFlzpTroSWRTEHPbFOYgw/flrbrqv/
llPYBUTDYXn7FQyAP5vnYQmxpBPgGXvb/CSEa46RuFfgNMIpi5vRfrWU0sGRIsQW9V05wwCZstyz
IAR+epXXe1/bANn5r0PqirvEFNuvOsJ4cmS3l16tmy3LoK/tcJ8aqUzvy3al/wRNRrwoS3B+038d
t+Kk/JBaL7CD9kYuUH6WAmSNUv1PZH82QXH0nWMxnlLzhCNgf6dQnr9QM8zscLmk8t7jkVX4wc1e
fwNLJF7th9Uq/mqm1gZ2TZ4ksQrnNamfAMeCMrR2zQMRvKtukS2d7vM2kSaHvKvSqG1GQsDxZ/d9
219gV5+Xic5yT0AFGG34qyOIzz5kcUVMIBEDqv+91SmRD+a/sIEBY7Rz/iG67ycYCZOuxvrHSL9i
dWQFn1jcbahwIiwUokwtnMeBDtXQ84H3X46rjjbXhi4fnWLTsuwqFnSAtkEQRyiXOdtIkucYLQ4n
xx+RapFurwePs8AM5/xrcE4QPyJl0YPbzmLzZNKisqlb69fyhG7puACTTH1eruvGJKMc5WiLEpZe
jMQktMJFksl1RKgb2ROk0553VUb6IWtHy3NUpeD5k6IKSSJ5+Tb9Q9vrcZgloN8gaxc0yyaWW4Iy
v87e/6cjEDaHCicif7dwQkJ4VWVlx5UTkgT+whupGLYcaGUbXrLilA+7ORqb/BADHOCLBcRS2y7F
o0jRK1sTUColieIyljioeib4jR3142Vk8XNgLKEP5Tz+GdoNYfl5s82+1laEKqWH7tqW+9t+EYYZ
I8VTpEAf1gDAL3yl8/G6dmdt45BFiNjyA7I103qNAObiAXopigN0PV7Il+X9cOqxVHiBCwpCc4Eo
f3Wc482TG4CvDUEiDLu9FE1BdsXA9v+Uwc1VCeOAREvRGC/JJeGusIMJamcpc47eYQwkQj/p6H+W
JC6CYLcHyn1bIASKy1ReDn3zlMV9BmI3oIGq/mOl
`protect end_protected
