-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SsbTXZiDTS8WKecB4gkGwDUQBWg69oM7lrrocSgZ066o5IvVgk+gFw8D2x2yqm+IpombXNSN2oaC
tFC0KzeEVg+3pbS9AqJBcP4BCBcZVKG8Rc++8Olmgh2givPA5PF2OQuhMPlxozlpnAp7LUXHu9y0
g4rlYxVtcgEm0ikLGEurmdZzAA5CkoIaHLrZCqpvP9gxhY8MyomOPDQX9C0xMHZVszbD+qZLLJ37
K7+XmcL2jJQgUzpV0PeurqJEro/HlBPF1owxVmuKpzYiWQtc2Uz8iz5H5oakRQOTVNP4abbM6X0n
xXumq1SUR5yJ1qTk3jE/DQDKDNLP/8ErZOZxKQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
kk7juljusN/jbS8M4hy6uq+cRexaMv3rmJLBuOHJi7KefIUCkIhfSf5K3rUFc/GpegxyqM4HtDii
RP+ozYmrvUBWbtvmsrPLP1cwGr6LTUF8HjGaBVtvDY+dnYWEmmj+QtdLFnjk0aQWsSxACpN5sE4m
qWsZ5aCv+MqFv1Hoaw7JqEi2lV3uWP/MFZqjTVvfyufE6JL03cpWPKoao2Vb8xISafxRPcdfQWRa
yQpGYfGeB69A54hKeUEhupkQEMe5NYR2uXlagBlmkWH1HybTAndtBFEPgg4huhgwDtCdHp+Yl3zS
YqEDJzWAI7Tyn9wUCW++/OE0W4MFWtOGZ5oWBv+zd6Nx2wcTXg0Xgshz4GAE/RoZHsrA76R99KQD
TeilvfmjXoc7itVqYjs+Zh4o1egKlJEjq0K6VUwW5UYUui1xbMB49gN2MjaddxnTRDn0SzfYT/uy
UppnNLBBocxZ2IEb5NHt+9CXM2tb5d9Npu8TByEdJggrugFE0+VboAlIOkQPBGyZB02fT2rK8IXI
4vqigQpA2MqSMjFh3ShHN+bpXvINLZ6tkumEDH9yIx4VlqIBNKNEhedRtE+pSVMvftrqCLtjzTiC
LQG++KCRtj4a7ntsZ4gZhTCot+c1nBR/BlIktMpqhgrzslI6/vOWys9cFEK64U38i8YXjED4hpsI
3+CnXhOXhMkHrRAbnywa4N+LSBtQ8adxw+ptGB97KxhVIaduj44yQJzkcht0+P4gSY6U4L/U6v8o
TwRshPXGRq+G7wS+ADffrnOEOxpPL2vgg0X5jSZUGWoPt9xnXUY29teYg9X8+uwy6pyLoy/Vsqpw
SnS3kjctA8gvN6P8YBnqoP+osX5l89H2D4M5yn4eOlsKitvJkusm2Wg4GSuQVvFljCE6nYFL4WJ6
k6/iPVtp4ELvKzIyQQ2lWr2eDw0xfFNdEnQZlg1w0ma+7P96CqjxmOEljvpbhKAM40fBZ2ED3x1x
0uXiTHoRIXKagP60kO05mrRWQizG4MVoz1Oj12CIselmndsWdurisUpfOyBH5WlWVKNCGm21/d++
INw3VOapMBqX4Ul4YAoTuN7y3q2ZdJcvCwISBt0S0/6hmK1LRQ3VubizyxhziZe5f9X/goqKDC7Z
FfJ/dy+qAiQblohkVTy46apC4n3o9PlSLnD8p9CGDccGRTA6MTWrgi8hWx9Jv/29bjffOLnRq6Je
CA1enfSo8sjyy4/pVnKZOlxqTzw6cMSZspBejexJJHkjLcl9h61pydgdzp+D6bKzAK/rl21UcN2l
Vuddz6mXVNmIyl4drkkqbFJEHehfy09Q/YRRScFoMY3BoibABjqhSrIaWXuEdAqZJKrGCr4xYuaU
o3g9zRXMB6jwlBYQliJHrq7SFrQIdQ0/vjRE4P7jCdqPLm+Azd4+4m52YH/1l9XB/n3Goy5GnBjt
9mi2clrUasqqdHeGZiaugjo3quPCWVcvdFG9t1nX+jBC0e8TFEmaJ+h6ZzbDt15UR4hbvCEVEVKw
KaWNGlqLf5PlQuY2ghLWtV8r4hS+f0GXeKehGD8xPIiLhQO+gizmaaAeXvSHjxGJtxtMCv9HT6uO
cvJIwrVvAYOq8Zf8YipOlNNjxouNqH9THnt6jtn1KOyVNvgJhACR3AgiYh2a7jW6/QFQfZWubCET
mATvgJ+aN5BCpazcgwhOrbpCsXtnvb2idk/pjeTatL0ktXbVNugDGEFd1iSBz8Oss4ovo9dqcGKY
REY29dm69m16qnFDXkrri6LJu/LrLMW3MVrJgyVIyhZiyc3s7s5ptlUiHYkTQTXnxbq/N9m1Sc0y
jWAwgCr0fV0U7Yo04iBjxZQk/Iy3m9bxZ+nL4gcVTiO+U889geU0zJAWU2loyiRYIM36bv7gwq60
BmEipaLaja13Q7DEZ9/7QidspHeYFQzkWLHZAiol6klovori17TnpoQIVgspAf9NL0QHx26wIiJ7
fAsLY2vtl/9h2Z+pC7q1A3kjf4SMqsPy66NPZq1L0BmKasPdE6Q7lWfnvH/RPzPLCg/5tTR64UOc
+oHfzInV1avKO7RK43XuZmUxSxwXtzqcivHtfps7dBoUU6lhBUN7yOmagFRrJoKyE3pm/z2Ff0t5
j/JmDgQRt8ZRJH37WBZc2+KiHa2AJ9oshxc2hiGUukl4EIAcRgmRP0c1tid6hdx1n5XRyzuucuXH
kNLTxLUTlap1dkaSXFC8USlGVdpj7c2bODzbZh9NIcVDjpuWj/JwfITAoBmVyJzRkZwjbhPHYl/I
N8wv86cWIrf2epxXm+JePFiTlt0qfgrlagQYn2rSr2wbczF9Ne+Wj6RCBpssnQz3oY8DD/+orjZn
FPHsBe5iA7KHkgcvYuuMGWi2R2jZXCBX0m+8W7pHSH6VKe2ph7czF6iDmiADQNJlYtdRlc1lqppS
xCVLh3CUYLQVGA8dM0ukuI99LRIOBO7UXq4Al3jn9u+l19BMa3s6YiBm/lyINgPTxHEWHYVr/CPq
rqpOXfeaB9vyrm8X1Tef+r3sBlk4QRdotzXfY136kNU6h7q87BLQ26klg2jKyNbRuP17s0N1nDqw
AuHi2Q2jSQGD1ph993COR6zjadSUiVERltMpfHTECO6Wg5KOoxqMNJHww4Y80C2tKnIT/dSXI4wG
7YVlVtNu5eksEgl1qmk/O740Svp+4L+mehmilEFy8dPc8tdTyQrmvM/eu6G5+CMOI/8L6LdSNWwE
+6TO42EosllgHtAKnmrSjIQ5aE0guucn9gR4Hiuv+OEACfwaj/mHZ+87GVmNTnJvMSWZfLkM2b6p
Mt8sOmHmnwd/wk31XiZHZP25Nyssy48TnHPAbzbLR8R2CFmW/FCFAM5GPcqDc9RAAxABmFEcp2t8
5TV6alI/ml9omDQUcRYJHPI/zjVGNwFJocFQpMwGWd1+aiE/H4/qoh0AtPddIJYPfE8Gp66Qo9HV
8CChOOLVtGhuAT4SJOnAzjYq+vumBbCood0rSfVwp7uqgFS/W9Gwwe9zweQphUiRnvySO7CXldNH
drGRHs3qDFM8zdfzoMOGyW9US6y7xwoJU4g/KaeB4pVIq7ekmMbqbBzjgVdpeoyx466T5JSw0lXJ
zZx2XJ15J6dSu3fQRcloakcLn5IkGIiNsw058bilx8SI6jCJwvTCzbmX5lsCZ9HdSt+vFx8bdNqq
vuykhIukR+HX11xUny36kMs8wSup7T2sQXU/zrk4nglRsZrbG/MhzjORVEu9DT64mQ6CgL9X4CAY
H2sZakUzEwZBOQYCAaELQ7mcuUHVscDm/ktOxiLx5lW+cazM9MmYODb/rMGppQusk+zeWSFvq3kp
r7PlNtRduL1n2UcYbxxbfJ1H+dx268lkHXD6Ein7m8n3GLl3ErG9w6yvt54sqN+V39YPLs5IJCLd
R/mQ0sUh3W002+6gcvY3ilwVDL6OYqZCPDvSZRUYj+EYttQL+HUcVq2EwG7jFBnf5sau45msOGYO
IsfdVkEYQRy3/cUI2YArkYpYXbW+4p1tl3Crz25PIFQcvGA3SPUBdGgECE0VCOy08j6fEnioxAOi
l95Qdizbmkt6zgnkALlRbZxEJLTZg07G30B0g/yuZZV2/CLPHVBDsfmKX3tyABQmQiXSx/0DNw7c
USxI51NCZOW2W1fxYojJ3hgbtReSVd83pFfGSpoQd25llcB/10NtLVJx8nSaVj/h/tA6PdqlTR6P
Dj/ZNNFnXSsfnDOs5ilizrGpcfV300z6nYBFJPuQHjAimPGUI4gclapDnkld2aAiFSJw4MQxq6Ym
/lpoI+XKrMRqLHtfZAr27uW9NXX/vGxnOfyIR7gl/gradQqDoxLVSnd2tf05PM47DGe/mel8bDrH
7Yrg6R/jpYaWYVL0H+b/QIMi7g4uY9UKAK5DNHPIiesYJrDvKf84lSoF2q/oy5lawMfTdnidtEfB
mkaD5JCE0av/MbZqp5qRILcYVvmGWMhf1W+OWtpd6MPlTE2JAbEfmgEPKrnSvI0uq4Lhaqqoik9p
Xum4gUuS//+m1lm+rqO99y5VSJ6+Fu86VMz+zUk379OKJCp9sw0iDHb5ihYZVKcWbK6ovInKJCd8
SoznmI90H12X0ng/QH4cYwZG1fJbkxEoYEZK2b4QcmWsPsdE9k58XTG93Hfh/lOOd4VpXD0fbDLq
+A01Se7greAr9NFvV6tpCwZ+pO6gXeHCT0gbTj7Xe+uyPMEJFsZc2hcivO6x5Qu+uljTEplGc84y
vjapDLZOAZe2tkRiu35xltEb/xCgkcEmbyDvktZM3oz+ULd0qOWmc1/KPTZkPfD3DiKVscXKHnCS
UDLApkwLQlwp0HAyDi+w6EFhS23K0VRAkrIxdWIpvQi8VIExT32RX8p1MY68FQzo3xbO+Xi+Smvy
jxs0LpecKQFGPRbQ+60KIG41l1ES8K4f8SsDcJvfwO+gv08K8SLVoYfjjqSIW3PNoehXMg4Z4e4h
y7M45tLRXwvAu/LljgVVBtt+LuBzjtUqd3EnBSUSBOC4ULmutE2+xOmHQD+qLqx7caHBDFwYW7GQ
l2ZVxqZd8aRdi2H2Ik8f6QFHEC8gcXvrmlx8/bNbK1koKkhe6ucMQQdcCnF+QODE8lIGaTW1YkxZ
J3+pxACVDHqQO4bRQKPqJtxDTKsPE4DMdYwOaaFbR4/TPDtgy+gzGOm+U6bW8y/o1uZbIHmSzPl+
drHiWcZrM8rA+s1llnZ1nqJDxeiZhtw3yL0NxW/dBhx4I5xCv2jXIU+jm5xrgldOjceKhOly6hv8
wkl4OY68HmJhvGyPrcWPEI9T33rw7t4xLE1CohMEDe23VkRtk9mLAerAzuDpY9WWJZXAPcIsYCym
2/KKkuTn88q8wb+zKSMwwVG8u/PAMeuWg89XN7GT6F1O6WTPCejcTVTZ/aBdWpcTHkpexnID2ixw
uunb6qWQJol/2xD+OLGd1dMe79Ml+N02OQImd3V/5o+knOVSohQ+Dg7FdIxzFa0Nel4E6mOvCfZT
83BQ+MoiCGAZwOOOlDxltwNZxc8R2Eu9Twf0eT17yxVmM16S2OvxYAwa7RZnU0ETxuH/NXh3HMpP
xrAvN+H8TBr80B9jUQxtaCWZ7IhlGQHMSdiV4icKXbVrfvqDdvOkRlXIzPcS9ytOXhv8Q4fQw2E9
JYjLRBlRqfmpka93uA9YDT2eZk85NP5cJeDV6BsCubFyKMvVf1xP5Uoeyq+bw/twNjdtWRAoozdp
Ce0Iz/gJ3DZtzwKa//1iZ/6s2LMorhuPb0RfEmvidEBdICFWMBWKR7DOspOecWGyKxtlIikB+ksO
oUa5BqWgHNgYrgDCoC2/9Cxe5qvkfjMhre8C3bQQ55DCLyJymQLQ8lbvXN8eYnRE036kWruAnYdG
aIs3MEmYUWTGF5U/yehxQL6S/r0oZUuoDtVIvpcC62TfkiiZRU0PYa7u1KkH1faoo0CUaPSEmJxw
lh+sgQF1ZrcvA1hcMHT47R1fqOrirCV7grofDER1gbTUw3zTH2aJNNT4KyW6sfIMT24OmrFrlX+u
cXSzKiqLUGH6Ux7/AR3CRrTz5eLbdmb2okD9nCw9iTpAYEDO1UC6z2KjVzU/Y+n7akJo8U5q807q
D7YzhkAAGQXz1ie7UuEveAUxyTi6idFmN2B5pkL8hhtYaSNifwAE6wKEb6exGn05EgjcbM8XuJDP
ri3opAfwILAeK74k2TMvJNeF/bOqI//K0svANIVSlE3DVbCMsOVy9P2UZNhjwimN6ByrM91O/fvW
gpL5c4Af1Ijl7O5Vo4DdekxMuT2gBAt0ZatDS9qARwSkLp4f7jyp2A/lPuwbkS5ISi8wcN+Mh22v
rQEGcjlIeSsRRQmWCEI37WAZAF2IFag6zM+HmS0x8KwPtZyW3jQVUhZPFgiJFv82sWEE2iVo+LIA
zg/7ub5HK5rareDOhwWkRrx6AM9Jg89l5/mw+Uyfsb24IXRuN0UOj0bGACxKvQO1s6FCyTlynean
O4qiaVcutD5PCAx1g/vYKibR0pnkMoMpcMTUlov2263dzh2h8bIFlx2S0q0qWb9bFapOWrBGbkWI
EdIZe9zaro8mVOdwYOnKouMl0QLS5mEST0dtKgLv1IKT/MIvuF9DYtWFBVBcYltNBNli6S+TLuDu
V6hV0eFhW6cPOZNpmEjOTR+IQB3VQtI8Z5kf7W9QUYa5s/cybd0h3WYxffA7U0dSVVyZ4Qqfj5vz
rq7yah+WDwCXefCHUeKfBLMUgTIXec+qNiw2/AwR1jG1ms1G79xMb6AAxtvXxmFv013R7ZYivzJ2
fj10GQLCXeWRmpL/56YFvnO0lBv7P8G1tpz2IvryCndVt3nyPOClZ3F7rbOPzZ5xo987WRDOO8kj
und9KBfBX3hXyjJm6pB4n7UhM6zFaKOWFd+Nh4X3zMbhYAINJsZ3GXuR+DFXkGP2X3tCu4hEkSta
mjnqkxW79nokU1dHmMeD1VqAFM9I6b7HBfHAphgphuNJrQznEGlSz6csEnMLyLHtd6ymt/IUWrtj
MLXr00XR2nCrwH1fZKYMXJdV+oJmA39W04l2iguUGp1nQ2wDCgD3SYbveTjomlZyc6jNdrz+WVlW
cnUH+/T1wUQCdUgGJlrQjfs0JqLPcGg/BQS5NRyfjyO7kzaZCT7fT5D8wlwpZISgWh84JR/wfzYa
+DCi7JA36Pxw/Np2Pet92T0oAAWtI+z6WkKmx+PwH5+RrSNJvY4MGHAv8MfYqFm0QZPt5Uo368EQ
K2POSxQaH1Sy/NxQyykjkJsqL0RUr/N/vqFdDAvfiwQbFPFOYyGmJt/7Xb4au4qxpop8zNHzX6/5
M1HWmL0AmuDQMN5yP/5NHw8d7o6SfmSzYG6iYz7Je8+9sZg+QjXvcK0GpiqW3qOdPIRZOc2TgG73
0ZkkUyHG+cQrdtJSEjQtqXQWx0XuEbifvBuI+sLmJJ6JJSGavzDOYTeFUJCLTtDg8GZSgK3I0muv
QEmTmGuQOIw7ACl2hsSLy3GWaCWjQ4Rs3AhREAqBa5a3Y/UmJpSyer0CXmm/3KHoVbrFZKN5AHH7
FHENAcxJRw3cLyk94k5uc4CKkhbV1Bcswqw4X0fOWznpeAXUwZYTr8hvdyE7jVATUwHzcQk2Zw/q
gToK+RxBBeait0tyAYShVXrunpV+7BHUvWzA+7Fcx4kvfi7pqJGEb8Sqcdp4OejgdqdIxyjmnzAm
7ARgaRarZRXhP3LA+WoSYBIpJng7jfnw6rRFfH7d61ivhAVqaE02cnQwhtf+ul8I4PezHS9dcDgL
SyfyONoUSTDAlF8lasMYLsFRY/lpPvm5u8GHluA1TCA6IPldHOWBeSagAig51a8EgTOvpCzzQ+Bq
XJK3uJYG3wVnXL4/4X4evCH7gXymxmKnN9BhVjwBYDznm2rsVcgE2t1OBnDug6WxjyBpSUjMAwO9
/RKqnWbkoQILsb+k3ndcX5duEq/XrPeFolZCpkyKw6FRq+FRd7uQz2owVO1dF1GwqcALF7AvYE+6
r4os4Gcqgxn1SEne7n838Dvj8M8NnCrdE0Y4KAZSbH0hgJJJegRNz+6RLdX5o7q52QM0XtFC5tN1
tKcq7ftYks1sDA37Ga7VwJ5itd6QHDIbNRqrWYkmzEhEY1vtdrqmA6ZrtE40scJVWVShWnepuqQu
uhNWuwqNL4fXg/4aJP3XXFBhOe0z6mNccyE1zApVMGzXiOFSPp2OAv7OTuOmF2CKS0OT0v8eB0CC
+gJbi7x6WeL2fwXH0q/CyE0QkLdRhWH0wK7y5w3EI0gINEPzwYlPtA5+hwdoOi2A60hjqpjn8BJA
wTAzzxl0aqFCGIfbQ+qtZf0kd0AofNe6KdB70ilneW/MJXvvcaUG5BA0Abf1u/fQ27DJW6JkCyCt
4JI9anDAvmqgH9GJI99CgF/pfdMCGVmggEgeF/UhfBXDkPj4YpHTj8VqwOq7bXa4nFCYX78Tc21Y
sCOErYHQ6Gg0Xh3IrjCDNui98ZZulGZ8dJzMzMZxK5JTmb4Rr/4seU8RijH1pr+zohAoJxQ5OgOB
zhg4lv1BkYD9Rgk62JirD77JHiPuQBOt1FCrelnphfhHF9CIEHJ+OHIiKz6l6rLfSzF7ha0Yb++/
a1+k9XlvEZ/xQSPfpvDGpk1CAAroOiJkXEkEqwNlhDYYwdYR0a27viVD6HcivOn9F5Gcwrna2ZFN
dIjSB2I8hXlkAD5VzD9quB4ImqnS3wMnriaT1OeVvre477dlWPuVZwrOYr1wLf6WtaqoEpc0e08i
wabW3f6ZYYF+pCZLaZrvlXYCT2cdoL2byPAKTMyBWLznp6Zwp8+oYvQQviP9Ai0BoFvNWnzlLdnO
65nczgfZpSSM8emPRfFZCAgx+/swYVBfeRO+u0zjqWG6Ba5F7OVOO2bnUdfuDleTYwtNygRIVj/S
1GGDWthiD8zvXdGVdlyFEFuhjXEE32SSza+Tcnr8YZP8+U7J8T7KpjDecpYN14H12xtQwH9qTjPR
acAoVP/6weerPPDtjmEuoH0FvDmP/VfAik9/hX39+GqxCanGjww2daSwjpMRiHE3PGzQ4cKcnVHL
ExnfdsyqVtTEtwy5O5e6tHva/EQPCIQByaJNAG/0EHDTqcqRE3EAyhWJH0goCmccodLsmAuzAqsk
BhdIVKJk3O3mJAjJ8YK470DGaKtymabDmWWiWPZQRkXWn4Cfgp5A5+BJtfZXDTd0RcAXU/Abh9hh
S1+CAoIlmYmMImH6+drvcg0dqE8daR8NiQYUG/VMUzUq5kxRlbmy/tZJhaxfUguGmQfUMlx9zzi8
0gLpeTOGpYsdlxzYaSWm6zC275cYVGtr+uGyY1lQ5Z0UkzEI57/a3g2PTHiYnhqLJ7aFuM62iXB8
CW7ZFki8pOIrVqFEpihovaXqsnImIGpHyzMJQTK2/fdnV745dYYztrlh1KFklr3A9RyBUj/Cprhq
WpT+GtQkqXU2gcJi6gnNommYDnGXiHKE4eAPMd+s8v758WdHbY1qMrddgEFbEKYrkH7xoSBla8l0
jNfPBjFHwpIjJeSbXiLU4COvammTujEK5LiDJOjEIux3MdD5BXeFORomhtgwqyrXuowlbRjwd/HY
CLts0Xo+W9nYSZ8mG3aHv2oiCL0t/S3sNkp4Wpx6i+SGwPsJhwt3J587WZE2dFmf6RiiDL3oJQNj
E4pu3Sn3Fh6sEgXMdrQGqGfGTrFYh34hlDShfDg0j52mj8kecFREblXGarqGToKKL9iL8tAD/rkX
tIy3RPmB6bvNd/o2Kl8sYkiQGQO14/5QmSCeuGV+b42wvQyxnSiPhcqqf7sB3AkC5Zhwwg2kJL4J
ehh3AOXCJWo6BFSl6KPk1jU3b41fjCq13bbKNYA8pyqJ0T7uCo+qWJnQwbu9EBKypjz7cVfsBKuS
sY97uHSD0HSfwtFOxFz43PIOlUQZEKHqdKVdpjhKe7ZDzR77LkQUMf5PT6KY4jqaX8TBT23JBgqY
j4OvxTpqek++jZlzTY7eyAv53CMVlzFAKsl7xgZgKyHV/eezS6hDGJGrWKwYr6rj5w8XE78rNpH7
or2VIqgW8/268Bo1RH5L/rwbk/SebIQsSZ53TeJL1UrFEvQk4lXg485pvZMpeJ36cukgsNJFAhaS
/XR5EYKoLDQphKNSWA779J27KfhiA40zCSsKOixKvPC2PPKXg5Mb7S1B+/3G/tM/pFQSJyA7tnXr
GFhQISNipt1iOsTbX+81hnrWS63cHq41EEvHsEoErEi3speflAVqUX7ZowpoaIq4W8vbeVudoX8h
uaW4m5x1QOhVD/XjHfuzkICBuesPd5MYYiUXatpqM7g1v3j3jz20OWaqGZvVwC5IL8gdQpWEjRm7
FeIH+dYYauurDIVtnhBTC89V7LWUUflvOpLQluJizrD0cwXmDZmEZYi0hB+NwJPNmDLyJBRj2dzO
2UgY1kw5pq4qctEzk5SGlnuUIvp6mujYb8pAfJ3PCJylkAyXz4MWMdSWI0BO5b6kNDrOnz1XrBLg
ic2FG+OrGLN2P2Y8xnjHIj82g4YwLLcguOi7ckAd+Ubylh3Q8bncZIIODhyWHVF+urV/UJ4H5x/P
euBPjiSRRGhSIkfKmIvbjHTVeLmUoW9vAhCJpN/g+Tl1Hh9HnCdh0G805HyYlaBeoPRPr5IimvT+
ucg/POXKrGEFlESq3LSFGtwYgv/57zwER0wd7yRX3FWVEiw7y98FijhjTyL67oHoAV1c6YzzFmT7
3IPPoNSI5DY6p2O5d4lNtpAG2kdlFk9PljUUAo6Ux+RG91kfNlD+VV+Jp1oRL04dqtjTZEd1gCUC
8G6ruwQq53Xghe+9+/YXyMPMeCL5sILpOKvvGJ1tA622nFM7g2JHddpuZqnUeoJYG8zlIom7FNVk
DbW3Vb7Q3GiFEMxEqVm/x04dBeg3OSijYrOa7kFgRkpZNKMjO57PqGS/3uyZTEpVBQYl6muts5dB
C5w+v7jz/cc9Pw+c336dprgIa5qSQ1fu+0y1Xu7aY7kjkyCW8z4U0QF0pBWVuF0JeF5fxGfLsaqw
r4vCTuScOTpeagsWVdrv11nNvAZugJ0NL5hb22OEUNwnVREuAXUiLL9V7lPokeLaFEzTyFagGXx8
4OlqL8ZUQdtnVj5I/WHkuTZM6dHK5XenBFa0EgystquH5c+EOwFy+cm1jt8Z3wgMOPZ7gYCD/73G
/wHt2vSznAIk+USNM4puTMesiUJymUkwkNEg8p2t9+ufDxqSxR5K1voREOVdaSte0Wb/ShPI3iN0
+WXnwstOrC0sSYKfC0YGls7N4VynnuQ/TyrOsZxq6As0pXbIi/K8NIOyzBSeBUBbNi8j78CP4BP5
8JxPXiLxHphAKW8ga4qXbVm+QxZ9qiPSdxcqA2eOS4h2WytLnKHwjU03+7GCAnPIhM2YxrCBo8ZH
wEViwa+6reNYtLBT8tPUXcivs4ujzY4hx7fgtyoZgBEdh2W+UoXxIf25AJqzYuDkUgIY4NLj23UL
cL0Pd1V5AKn6n732dBrr52gGZLrTivyooiu1HqRKnmep/MCh+cpseZnZd6GIeHQRZI02UGN+jSun
p6E3p/v+xD3Xjk5kzlSi2jX6ITAM5AxBbNERJBsw+WN0I+BVXcAf+Fqe6Bl5QnBIHwwX3zowoEg5
7eEksvFoRLBqOiZyCKHUY9K7YkBC+CBbiHC32BzbmSu6SzI5v6YvJsM7zFKv4lOKwk0RKXuoMJaE
oLLHpHH62ltQ/862afPeSUP8hh+3ul1XMGswdbkLCvdIMTyvpH/v6bhT9usR7s01hVfJNJLzzlNA
h9ozHAoQuMbxiPdjFNANqDh05XX8xrOC1msCCHrKT/lsIq8QXnb8RCSbL1Qcr1KaJNPnRPtjalKu
/ApZkvMfQGaCM3l50X+2fBHmoy7HxY1yIIv22A87h3IQM4XjZecIhRkH89gI04U2cPGVcDRvolc7
zLviMLOxTDv/EAYneJsl6leGHvI3dB1JBitDZ00Jiyol85XShKZtXdG3Rjn8MbjegAYD7HDIIBiC
w2drYhgYfn6vU82CHrL18JbbwbjDGYUTt7I5fJaj2uBeNKjbJ0tGr0/3CpYseWQ5Mkjpx/iHDBhf
th2TexOChHQS5y2AnGeQc7/vvSrtc9kE5a9fSnEkR9CIE/mwESE5ZHr54lKFW/PcNZhj9wq+wQ1X
CC/ATHLdBoruBwMvsendERBwvHKXlpnbC9FLTSoBMqJbdG6+aBx4CAZaFpq++Muz7Z5R5VRqVI2H
+zAUZeycX95BPwTytb/SiEs31YjdM+1Fem3+STJESmHi20ZgFuLbIlYG7BXsVwPHlZzGokYsBYRG
wAfKwgkI8dGkTTh4B811ECeU9AkloWYjCrC/YwKTeWSaVdSk677hpgeNCr6arMTreztAKljj6pr8
zc9+UVyjEGjJni3tXIvEeKUKc7wb1uj7S3ZI5dVCOotTxx3CwnHTAQCrezaROtoh/bpAY5dFZ1z/
t8eNvmnf0/Jt6eiKh9xtFCKPR3G37a/YsAfiJ666NiMs8oKFTsFw8VfOVWFwqI4tkbgrrbAWATvK
e+ptQR4Rr6A93tkqYOwypsMIaB+VsIRCLyn6VUcPfI0SY3nmca37rjQoEUt2yhlO7cSEa7Nct2aK
pYXY6+jFqYOlSiaFGt1u2MFrFg4g0Iv1Ng4X6oMdKovTGx2eqxQLzR6dWoVKq3rgLA8ldk5deVnN
n8WgSfJWnVVNZXkBS7PwFKiWMJMo1OJXqXOoqlHsRZO6e4FHDWgGnAd9R7YrO3x1wmeCiK5sAfWH
mDV3LAfu3Ev7CZCaV8rQBaHdDRAWpq1yVJeqTXR8LXseDAgw1T7m4kYSRwOraZPH+CnCspHSYv/p
TuB/3b3UF7Jqd1ooIygxfiYJsbd0HsPI+ro2AZIZpsmW4B5UDuAJbkB619DRpXtdw1fPUO9CqsuZ
LoAc1sxvbqfy2DcOlQ57ZOYuHWJ2Pm5tjHqT4KgESip3B8y+caHL7AsgjThO8M/rY9wt9rPTxtlR
02IrWTpiHy7rMoFNqU6Ios85aUN9EHeJKUueyb9H06ckcHcw/VYgctdtNsLdcvit8TWVTprxbHW/
WIWXZ7+qi3TGczxGrbG5CsxU89eOGnirnUS0usJVI3DlVXU0WNzMj84O2m19oobw0+1mZQ6XAqHc
Cx4or+/qKqmDWcTwSTHM8wqLyuOZkzcRSLoNej7f9APuO0s2QZ52qsQMChIKdpqPLj/nbwIwx0uD
Pnp9PlvLG0F2KWanzwPRdz5awzzhU+rcxkgiIygpTOB+y3Fb1d66+ttWCN2EheWJOO26JZ+PJRfZ
IJqiB4+u0QTUWvfT2EwteMCOYFYgRDjhQlqFS1FkefEEMTWOqZpjA8NcY+pDlrXqrEvCT/D79hNe
zknR3aMm5WodsVzO/Zqn3udknYqoDLSwwb/G3RXqGnf/OXbnEuBSIiSSCLGg33LjJZM+XQh+5mf5
Wpw9f5h/s1zukvUdGtweZ2ejQMGMO+f8ASlYG2J7DnqEtdaEb0Q9q/3JvqocQT3cmOIx8ChrEi9J
zCiBONVAE/oRWRpKO8TL3I7+ANJIs/eDTMsqyqmIrYYJ6rgiNXMMiUke3stKahyGW68b9m7p4H7w
ifU9Lkp1aCFFp42lVGzk4m1OqAAPVXT400cRbDS2lkM7KU9YFmiirTdOn+KPhggvO1e6gtiMQFal
FuP6haXMlu4q63E9t5WvtdQ93xZpZ7ikjp6jKq8zL8QVpqIrnlPS3GaKZ5eyAUYVqnTrcLufW0lr
Vk59Qeiggl4RV6O6p34JjNAdkSO+99Ta6Aw0saTq//PzZ/pdRXe/6ympb38wq5vTPzeGX86DME/H
d4kq1MV4ZRWLABc8zgTGfbCz7p+m93QvkADSsZQS1YC0zjXFtir62vr7KJOqEp+kT65dUjd0bFnb
kAOcj0rpQBxnaP8ylOJfrshF6mi72SrRY0RE98a//d0YBf/8gm7eCH9ym4LYnOFZ52mraLfruvQR
sOJ5GvV4rY3xSYRfbYE6QexD0vZS724tV2Ud0Z6L3l6mpqkmK0zTmeSmVRMIX3JI6Z6zarBET59i
sugotbWfSdqzsOWKgKHGCmayGDtDqiP0mSwdqpFPkrI+pabSOHuGcTdirQwuRjZGNrobkyjIkTRJ
zdPHgjxCoxuROHhfRcCZPgDMWKyPGVpG0LF/art+bLwO/sQFvbj2YNBvdLGv5ZE4l4LuAX0M6oJq
D1Ba5xrKLRTPUNcqVfvS4jj9XUaCjSPxmVsQeaKvV/y5EQ6HIyf5aIp3HChZ7ffKHFgYXwZJpyGF
ULOLyqhNx6xwK7P6FSDomkLFiA2R5DanDLqPB7MPl5mi7vXiJ3r9wLr6s0SO2Gjli7OQg9646WKk
VX48ABhp8dT9OhHDstRBXpzZAD4NEohHXwjD66czpJulbydNDAdikMfwo7A0mKAMNJUgHCyBX3Mk
AUkaMlWpQS6VQ8reMM313ZHxzK5UEQsIpLmQEamcNzSRZHpKQpNyO3VC9X0ygsKrxFC0W5PneUh5
0/G1ljMckSMSEW9jP8kG3iTdWkn0LC2o9VDPU7JLQoFC7vHO8kbybvQPxFE6V1riZe07hTcc64lu
pC84RxAj81UjD8Gkg9D/K72cwDMyaHh0g9EQAbQrlsopRfT0xBB2n6Pt3fbpynGeoq7sboYag+5B
3kbIdnqh9fRsgSz6RskpUNBsgz8g3f+PnUTQdNL+v11XS7OFD5DbWaYUq7KIc2GEVoQDgfM8e3Wo
F2DIJwrY7VioApAFc2JvPqUDxQhZGj0/7CrW1vxBhffwfOCqc7n6UnDlY5A6PebLC8cTHIdMJJdN
SjDpjVHv2LxVGcC2sMImksC9YXj+/Xr+p1LI6tfN5NX9nlu0VSG2acYbxqsrN19lKZzGuD64qqXv
RDpjynU4ZVghV+MHEbHYjt7Kz7RNXyMkm6UkT2yLY+tOI+FgCCAr8FgVYbE8sfRlw1g080R01o2v
NFHN54iwEzF+Gymyr0429wPS8OUoQnE701mtGc+KEfjHmnfM+3Ks7Oo/adi0QM8NUs/ITB+RymFs
ER2qyTnWFzcx05J9Omgf61E6IyR7wAligtz/m1NiGBcQXeztSw795QrGTm/ntnzIKey1Zs/9pLsc
dT9NWDFpyPKX6KKGb+4euPY0mlbzFdekZXjHdk41xox5Y1KDp9UQeGkfm/QwAmC19Kfg+/3mVmOk
xjj0Uy6xtX6msuo0FoGWeBqbMJcUXGAmVIqAdhstcFf5KbZkObhfwsrgJxnmYHvZxj4wy6IKytba
bMNqlEZbXIz9HguZPSvVr1ImxiZuM1kGK+K+FBZg/4ujNBRCLLn+CDoZFO+T+n8rmZuDZgidFpBw
XGuKFnZolTMaY/FXTzl1oD/X2nxsN4pq0PJjr5MPyn8+d+UpHjgDIyXfGXy7YTUOWMjE5h9TtoGF
lTYh+qaWYpMLpsczXWkUAkgcxVuNDdQyu4/ThG2044QerVC3AH8AIlWO2KXU57qMBm5U6avVSjyY
DTILbkrMrHwOfrx5PWFVCUvtCQKrOrjaYeKB7E/nj/sqcQ/CzQBG8U8/BcJfQ9wLoxwvvRzhJsjw
aGodT8/C0OIk2Ccn0pKnz5ieOidZMTcvFgkBXD2T9EUH8yW3R5PKlqG6mk1m8eaPrZVRRN9/d5S0
aSlxUYZ7nwWChgpfgwmopETB67iFIcPl0Hk6U5OhQv4JHmrWLl/5BklTZp/SwVoeP1OmR+Tn9z9o
ALWc3uq3voFg3IP+3Cl2Rn90JwZFBflFL5b9rLkThP/+ant7+VmpDr+XyLj39m4Xj3Ja8kqj4kPg
D9btMb7bKwukHUGpsixP5nV8yRf6PRZ/NJZoBA57Ib8IuxkfKkm9/W1CbuChAS/ih7W6gRCZVECW
QGkw4mXwiQQLi8FnJ68+j/VO48TsF4m+v58USzL9YchwLe8gtPQTsbrwVFR5GZ0H75ZQz0BiMUn+
e46irdTLq7SwLzZeL0UNxv/ycfCeUypYWNov1zlV36DORktoqz58D3pZ0T8IUu63Z6pc6+LBaj4g
Mpvp8Dfct3UXGGO6Gk/fDJeubm58/nVL+mPSUmBruIg7rOWEsRhQ7+zdkJn6eiahQSD8y99BHjpp
+w0HYPs+V85Fq//9PdacxqzMhuWZL+A70hAK26S9HS8zuoUBn+vBRKo0zyDkk4zUebIOvCCxjpmA
y6LL12DuqxrCcAIdKoY3FRBa4ywBXD3sPbw2+xr/duro6cHjnZArCcY2iUw3mHkVuMrXCchglA7j
X0mZKP9uk9jIgQPUDU5KwE+mvghdDq8e4bo6Qp9CZ5/Ro+1Jgdkr4Df5yTkJ2YKyZPBKEStsEC3R
RrfnjS0eWN77R0z0kzbByZahVwLRVVwQoUTKsWNyOye+XmF46g4a++tfRMQ15mCNzPeSz1FICMVK
zREZ/E8tgnJnW5xPV0T6i//0oZVFAJ8orgK7aZCVAwaKGLzvsO7oXaR5qY30d/m5xmPvgU/YQ8Qq
+QOt7r6xEMU8KymM0Q78W1Fk/A97GMYqjskMARATz9Xmtar9BZsM2KQh8ahVuNC10PmitzW4r7YD
Lmt0qHMI8vGo5oaFcjPt84iXh+Yh8NeIGpG99I6XTnaT9DDmiU1rhZUDcm+mf1cRTn7Vn+3+NjLS
4VoGm407LxGpMufQZoaDVq0uIoQBrXKxjovFVujMb7mYJIEfTI3yNVX/FcOvJdcWkAhOj5Q924by
FseE5ESJSuCjGFd9p9lwDmKvSRuFTPcALOrT7cpF1rTzSJlw3Y2JHKygc/yYAx2EcwPPZgfFi+J8
l1gIYhS6EoHRVNEbeGhd51UbOnRlVh2k58utnRklReNJuQa9DeSKcB31sOGwA6IzeT4dXk2kFzmJ
P9RwbyMX1rnxeW+2cLoLzJIBAvkwmpZFVL+0ML+s7CvJ5b5fpkWGyn9jAAb39/l0ROfazSK57soi
aFYZ0Ue9JxpIoSUY2T8oOblEo8DtDeaNmqFUUAo61ih/CdGO/QTzG2DE6tZH6XkWe1bfPYYUWV+R
BVrwi+e7tvZR8vinBZFTJUqRNvnmiGbHORHU/ZsE9XsFXfyViXIA6kbE1PpEHPfpUA58JiVTwSQd
8kHakIdKXcomkwIlCjNnidd5IVXxdSfLMz3GvJm/3OufTPWGf5XTDKaFbj3hcpYMR20MvQUTVcg6
zkAvvjd3MbJbrsypx9uVFV7vtZsh7UxaEfUjKtU4kAQVnh9Uh1duDH0sgjB8rkNkIRX4WYIJNqWp
SiAYmBxIHZBVSPMi4inlpK6yzwJu8p7yHY9H0dRgMVwR2Hqa2fS140N2fzecZ7L3OkWbqBTI3twZ
mEi9p+Es3gnOuJeA2n5H9p9odB9mHyo9R3/gtMDJD7myVFcZvp/850OljmmN889iNHlq2HxiRxBJ
Baa2N59srNRLOuKJmFZgYsm0Aiiuc/EpmjWXVGgck0vtn9Ka+y4d7Rsu7yuk5l2eUpRm3wKWSFcG
0+hQPcnimPup8JhbKU4FHIiN3WqqggqrPGtdhk/FyrnkOUBj89NWi+BUV7IEzSEqkQsBheufGrtE
ocYnJmA5m+6ALllHtm39mnBd07vf42QmAYCUJhZ8sHxzNlqJDcUTTxnKnxA6fNLZyjGm3HGWpPDl
1rj09X9yhgHSFiX82LGYdVUbycGDskzd9kkyRqzvxZAecXHp0oLUeCpAU44p9iLFJtoJ1GOSsaEH
9vpOT3V314+5rogIosHjanagTCaUYxoKNYazp1KmC89Rig4dZX+V/+lkwxKHaEk349N+gZpFavRW
5PaykupMrGGleSpxR1o+IiM0fgXUV8o0OeouxduPA9RWVBrJUIOU9ulyYHXeL8k6C+rmsiD7g4ue
VOskHyI6DlNhhTCSCNB+7AyMY5G0z2Ht4wBkzkp2phizY5fcnfN00FHI1bhOlAsZz/7Jz2lSlYrF
EB3JWwodHfFteNIQ2Je+Knh3bfk6ZozS+7tK38nm8qZzjwtHSV1VuWnxq+LqCxdX/vXFt6B9UcHG
VHxNQIv/59mvpNnruVrvudXNzO/Ip54zjaAcej4M1ia/knmw+Kq9+/600aNBZvZNoTDrzoZpNy+h
hVYVXcrXJ0hLb0RPAZTVKUiDx7M0eWxY4W1kAMQExcnmxnxfQAo+JoRaRwpVxdUCWXieDI5QT/Yk
Kc+Ol6TPYdqhtTA+1GyFs+nOfc+nLBGzq9U/wsp+SYuZMl8TnbxyB0aJe5SWSnysglxvDVvmDcYD
c2Gf2X8ujrWRNECmODQDYGPSuMaA10Z1aJBxXbiZAG6uKCjwD2mBrhWb/5Q9InOZnSCU46+P0H1F
Fnm52RbnOvf8QTkJZOYPJlsWfnlCcKGGLkWFIupouvLN4l24hS+fg4LihPjE4FPUUkcMz6ShEG4O
8ABCb+3n8k9l4gK4JtaqSJaPT5NU8SDYpIvZjzQkm7f5kt7/biwIX/daCA+Z+ed6+s0pvzcvuqSn
cbGPZkkfrgCtzE+X1CinluvV5X3CaX1NID2Ya7Y6Qq9Hhc5evWKSiTfEAmj+Nw5raTeddjn3YrvE
A+4FadiOwaZ3x5pXl+M/dEF59cKgZwjjoNYJQvttVGzJNPc7Zy3wpbkkBYwQkXTHyi1V14okyJdu
uO44qxjsXxTVAXFxTOHWat3rR9kvlDCzy9kKFy502d9/+S/JNcUi4oUO/xzGhU/WjezBA4Ur9Xg4
o2/BmLYc26D1n0SutkllOUvaHnkkbeMLbsuMM+Vlk7GnJIwvjS/elCuK0tRJJ5iWObweW4pkXoZf
rgB6zmb9lqUPL7rzX1N1pWv7KASXQDjEzVZLx0gWA1zcZJhT7UA17s+0yhgF5c4y6HN7UK7DTvPa
gDvlekNQDqU04ZkkICQ9CtgCj3+L3F5LpN5s8oYanixdMoyRgMzDb7aERQvA+bATcyaJTc7Bbfj4
CnMjcsUyrpZ2OrtOXxIXuYk55x/bW+md0Bi2dq0FeONjGvb9vhhgE173cnqdEFQCuojOGMvpuOJh
aEItPA9NWbql+oJuOQ4LblvSYnW3WXxnCEW+YQqWt+VjZZBCalPwnhLFCLeoM1D4igMhTm9gVt0d
LntLk7PstkhjcvsXhEJo45u6n5yrEgKPnmHDadcgScvHV+L4geZtGC0gYURwHUN8+tV3EYoGIZXF
qKaJ5LILkSpl/kxmvFyIDVD77KN5UXpUKk2w4A168J0H6AApVOvAc1BxEtoXBgX2hP4ifTpAIWQc
vByPOkr6+IIL/AKqEO35t03sRj3FK8ENYFUKSoX0D5/wXtK2qzdfcCGJgUUnSQ+7F7jj6gRTAlD+
8I06XhuQRRhwHQfIwn+zY9lUPJIS4/JSJRDCgKn9mgcNZMm5LmtMy0SkW4Fk+NrtPYSnBPoff3Op
YOX2sd8i2mA69LkLEcTUa+YXoR4PJZ9Fvw3OczIVFUPOHmMVDFA6Qq/6rprQF1YrCl30vJq23KB7
J1xbpe98pB2N/muiVwkaZIP/OZBN9POWoyoSF/oxIwKyQJnM8aObGkXcfMT0AL7aMkGhuy/NZFC1
SyvT/42ivonNh8h7Aa6o1ZOhsh/G7b/AC7ZhQx0qy7JzKmiDjoULUVYCiCU0NTOPFZ0GnCVGSmnS
yvKM7CNid6oSmZdsGVQqOnip70U9zx1JYFI6e2alYzhQ4svX+6wVLPZIgVhZXFzprErdZyW34/fG
CgtRWMLm45xx28y39dx/MYyOZ18Bc9tI72DrgMc6i/lzGog3HpCJrIUefur6FR3WdyUGwNxpLjTU
c4GBO9tM4cI9Q5ie5RVw/wXFgyMSozttfG7DBepwYfCuED4sPF73vTId+etiOKqbYtybkN2lwraW
ZAyZdFqYywVfrCejXX/k2Lnj6GazDi6ME65zHHYcD6gcTd1ycqv7g1IxC4QrrsM4abnf9EBxKA50
GmJNLZvo1Zijyhf3drPxD0uw65HO5xZPdynk/upXSZo+9mNck+IMYSpwTprGSR82DQGwJM6iwX35
ifGMSh3/9/w6xZChpiFRo2CoIkXUc1+rPucdNo0RLdUA+k2UmTqk7q9HL20LDCgPAv1LaWVp4XlG
c/nT9iUgbo13CnG0ybcPH2RKsOny7kEh3zv8N/ripdLZC7RE6GD7uPdDxFQ6Devb0W3lywMfpwxA
eCbJas0L7pDahGhxcS1sCz3C9KWBqsETP6qW83lDW2l7/b1QiGlnn/AgoZlAoJvIDscUtUyh+ju1
uy3HrG/P4hGkwvcUOuRloOdWff9ybMjD9EWBCi7h2ssYyR2Q0pbnwkEJsi0mFfP4DHXFL+eg3hpm
ldlXF4zB/DgHowsvgMS5G+00C14687fjGG+KcwFG6T3k4f6kabdtQdRb3oyw8vfjUeiRhS47Hnm2
nPkcZnZilm7Mb7bRGqgiZTVZt5eCWlaOHBvNAyY4NlW2Iy2xYJ0SwR2yv31tw35Cjk50B/vT+NPp
ywSQ+7Rb7mgMhpzm2EyyxQXJy2nbORYoPatnMebW79F/UIUqhFxNNjg63lmADs6fxWTOj++ZOh4p
CvfRj4nsPRJFbfyOqxtG0++YWPrk95G1b6QtHCH8r4I615fpPSEEavNyf56L92NUEdk9ClzDwGml
2MFpgfKz/04C9unztQMbrKlhwmLMgvHLsyyqDVbF9Dc23xRadFlXfYIafWIwjPqRZzliCO51chc/
sj4RYz0hxqukSdBRDbf+JTjTRplPpIq3PvxhjNeRxOJa75hWOzsUAyLF8+4FX9gqV4+wDA3jb6bs
Vor/cOco4MRK3ltwu6YhQXwDyDuMdqYJzyKI4jwyfNz5oXH1IGwj3TueI4WggKib45QIx+p1dQhk
fjf36IUd3LGgJiQu4vXYLQIU+vB9YoY/smPf1PIuCCoemDt/qp486C5tQ6ouNPKy+BzOJ3Gv36BG
fuCHvYC1nQArr1hU80x+7pqhJUUS41X4MWvwptgpMsBnrCmxtI/f3JUWpHeQcfnTLJFaz0F9j5ml
1jisR5hzHCxePAKQXz1DsycGybLkCI67uTGMAK3KjPbOMG1QV+2CcouSttYlvp/ukUtm3QndFcWO
7UA7Jn+28mNFGsOgy1twj+meJ1dDxU2v7DPSoFRypN5qgH6afFP0+jbweAON8FfkdgG8tMnT8/47
KAM1bFRiiSrFXZk+kKV2Z9Fu22XPUSkR93GNn6Azc4Btg9oekDNtk/sy6sh1TY8bH5gY7DpxgCN4
QJdV+496zzox7neRvQiAvD2J8ag5XeiSRTUA7MPx9/Iak25/3n6og4mF3Za1j3+X3GZa8D4uiMTz
PJwkFZmiiOycjmgMqqKnF3DCYRSOwe2IlnQhpezSUOIki10EmQlXv7iLjAnN/s9j8irYiXRhaaWj
NTxDLfnUdHSoloRJgiXV6pBkDghgPxxmvWBlzYzHIEv3gCUQHz+qsIpoxetWmfGqziruLGpIfNGm
5w/9SQ76UzOAzHYVpRCvlWpNZoJcbJovUnvVmUzINJFPnxQNpXQQbGYlbBAz01KMge43tC99PaW3
gbDcvQ3JXAXzCcD0x70tQpIqBfagxRZwEMW7ZXliVT4wf794hIFqCsQnb7tF6oLnW57qzig4b2N5
zdXZ318CewUabNAATti1OSJISenL3JYu53zLGlEP/9g9ZeG2G65BIHQAM8brb+ESe0AYGBsQPFXO
hTObJyFf41beIac5jXfjsh1rPVKDpGQ0Lqq+q1YBV4zN6TM5P9MNlI068oszoINYCHFYEl29zkHu
6GYBdjnCIybOAELwMX508+kTmbXH0KXlwHxnsTTtMMVpoNjKvZX5ucvHqq+Jt9Ivnrp/iy5+BM0R
Zm2uiewCNBl7vJWnKe598UTgTHrtjZ7XsA00jusQmbi//P/nPMOSG1xpgX/ZKUMJsgw+fYCIfd6r
uvkw8HcIoc0kxxWi7pY7fZYxkTT5o7dDW4boXmBP019GKWJsab6mGPvq1Ci6/RbWGqLfDNCUoArd
rua5ARvrNxt7Thyj7k6G5OYNb1RDlN3LW/rxe59honHhJOy7cqMDaRwwzWViSQbvNLArz7f0RKAy
5M5aIwJmpRAHlx2lIvqYlWgt8yxRSLEWXII7hvDo9Ucq1gUBj6Cm23uKZK7a3mmqvk0YL51CR5XQ
UCnAWWGRIhsP8YeqprV1UoFF5O2ru3Fh/RAQ1Fx4J9AHqbgEOzXmPrRsnFuV+JXuZsMNoDnlBTG3
xDwkFZ1dYOCe1ZSji208zfNJNHbGvCv0DgpvC159z4ztHooq2USLe63aVeD3g+HdiV8zHZXtAIe9
nait9/ypmD/wHNJjf1Wznsc6kRB9B21oGN9PttE8/guxazCLfOru+7l0l6oN79UAxRm4axreMyh7
eUcUHD9S+cC7SGCVtHridr8P2/VH/lO+pYrhZyyNJd/NAeZkGylsYqsTE81AAcm3O4wPIJMBEWKO
Rw3Pn2jrJXkef/M6mSwOt7tKibJsHJFNd3/7NORppKe19OuBtbh7GDTi/8LvxHdEZoYVNWETWe5o
b4u5bPX+fCcwkgHkSfAhpIbvqqdglRQwjZKXm9wZxBGEQGepxKqLxUDG2XgtsoP5xfET5QNxsebD
DuseRAO8NAD0nHJeAPOuSr2Iwt55HOcZVVLyeZPjx1tw1V+F31Ox45LHTGM/OpOsIccngrqREg1w
DEsJHlsahJ8pIyowwnDjuIjxZyCwRQMGClltzBYGaHJvEN/DfrkxpkAHgZjgzohOcCru+QKhyx0c
+hrdOEjmcMPYxS5d5+79ZBnHVmaU73cI0onImeyBLx+7HR8LvmHeOqgUW8V+Qmk/6TdABAVNT44R
gLgGgWNbtyId5LXRPvWCDzVDMF2ZaAMQo5FK6xiIj06ggfhbSyOSRdLftx0zkM5xUC7bBo8jfCjG
cIRlGOQ6wa8aPTKLIMBp8bun4xDApiesZ4q5XmNFQbk3eFWwDfTM18JWq76hxCzCg0CLeF0cZ2Yi
9nFJ5eGD8Jn66R3kguV37pTTXo+OM2KpMCv/WCPic4Ks9XX9EjkdkKMOzoyU8PteQI2Q4S+fF+bg
TA6fm45JaTrBzI0KYdn7Nb5pZ/poC2MMsMQ77Yo4M4JZn1chreeUCkipsPl++b2nzAwOefjII+Tm
w1SMnpvUK4ZofZRKb6BC+j2S5zfQto8lR+GGbvIMudcSOcYyLm2DyIySkY7moldMUDxI0C1KDdGA
AE+Ty9jPqFIfzuSQYsl2KR/D5O/jZUgzkRMNgrAkGrwbjEDIlZG0Qtb+LVH5P3q0bAWqVLjLIQFG
SjO9QBXj2dOREqTYwX+ETOkhIV49rqOtkrn9xTgQsisIqzwcQhE193hy/h/UDtsbrjPXbvfiAhzO
35nos4BcO4AYxKV7tMnzoeRuJ/KgSzr4npvo2DBo64j5YWNuvpRdPla+yHfLZpl9rW2FXuwquGb0
WDFOD8Xg0TDjcB4M1b/eaUxpD/EZ8S4QD2o6Tb7AYfTobfZgd3BZe4JbUegwFW6Ry2RBD0j5V4Hl
m9VZhO8Lnyl8rpyhuNJ1SS30Ao3BVv3ANA0f6DQkCXpuq0dvQeEZqlxKc+P2IVjXkxpw7v1rkzVv
zOIVgQPIixaG+ScAhwC8yxHCwBCAbgXIIsLGdid/PaKULkqS77hHhUZhWTIvHv2vik9isvRsW3Ld
qmx2qcih7CTXJhBTbeu12PkWFHabWlTRaqjBDoMUOw1Co5akpgC5DmQug+q4hZATFKWCy5sOqVBc
fsS+tuVtNhhX/OAHS7lfo+ZgxONFCBHIVTWO3L05BhVyUfUr4asSZ0efNI4ZzaJ9sQzYIp1TLQZk
u5CY7JB4d3fI3MPFAbB6oU486l+CSO78XR2LuPaJysi5pse1hYHAFSckDDabIw0nBA4TDrIko6l0
Xsmf+mSbby6mA8lKHpZQHeduy7pX5x3iT5ZV/Ib+e7M9LSLSmYZVZUpnDVBd492B3HiDflJSGMK+
6DjI6Rx41PEhq41lodgFeYpzOjOEaV1gRPPgy5Owos7eKYkDU+Ex+6bMo9smjY1p4oBmKzPqroo4
G6ICT99HkTgqO0abBhHWP/VGcrmETbHSw8jBxKivQFNHjDvZTGulzozKcG7hsaRNtNs++2FNTKOB
UsYACOQ9GSBZj7S+wMWQF2w/k91J5XwXDBDePtTExUzxuUyqwc7rrJw4TuvHR93R20tRkCChluD1
Et6KdVR67SgjjM+dGaWL/310D4zBC3U1gieLJe9jd/aYErR9AuPgK6v9dGJFZsi0Jns93qNLNMeG
uC2pgB3mJVVPRVFob67s+hTLoC9kHSTEIe1DH3xirnbOXtOJvrfY9VD+s0NJ58aAY4o8CWVaVgCL
NAKI/kh1wEnSp9m4pYB+Nftq4kvLAquU0Vv74RAwsB6Kl68mEB42GEjzwqoIiaEthSBozeJhPQsR
XAhs7tYmUqmutISSSXZtu4iHdq7cnU4+9IrOtYHNaCPO1vQCeQ2k/bJhplaETGZ+LGuTXIzX0EcY
U4LHqnfrhoxPubYVPxWrnjNbTODk9Z6mT0ftN0qcvKK0F4I8LLnRbVpHO7yfSAYL9WrXeZGV5ag0
jS645ifji8lpUNJFLPvt3Cy5BLXECZ1wyFq340kmqYCkcSALvvq711pkFR4RXsEbA2plXoWgLn3O
LVbVEtk4gbSOfXnYrPTM8jyn903z4z0bMLgoEzkCrIZES+jAmH+mb33nxNXO+YzMQzQONm6RzUqh
+NxqNCd0SF1VOOZfEiZa6eTRpy03kVscnrV3YHBO1jwq2QJzFw1U8jb4/j6aBT+IE2NQNjDUssoA
1jzI9f6hpxWceirszzouKIuU2Kd07qIYv3rCTOvDbY8ZQKx7CnECAs2cReM7LFi1xL0XP+ltz9Ja
4TxJYH8GHV0GYBDW7YTVirlhgwR7W70she5ufMvcJV1ZbUbiaRBVxsNgxGR8qCuzBFOpwgia5Pb0
mKd21s6OmmBA/HmwhDyfQtnqpYK/F43qfrzkTrD8rPF1nOhjRAHsUsfAcUOqVWZ4gMGm1QcI/02W
7w5ACy0n0EMlCZWu0h/7uY7XXbgtF4wDlW78h/uPWdWbdA9bW8LR5lW1qChn/9vvTq/PCwVx4NW4
NS+axDgl3bhhlCkwy5HGu/3kvojrX342mLGwXvfcWyGZFTXhuKrbPTGuSaK5t8u0ae8I6N5qu7us
jJ6YSDHlmHMQa0c+KOCMQy8IA4ORdEt5Qeo9du3jWJ/Ngr6h5X+M+U5vvuYtyWa+eZABN7aqOGyu
oIIYvP0IL1ZPOUfLAv+uJY/Vuai6ZJyKYTt/RelDJXgKlBhFpijGCiAA0txemR3WibBcb0WJI9il
K9mPwDy1GgZO6X2VLGvZPK2jnYb0369dv2igNNug7hPLkmBl7+XIYuwY90894gEor8sxzbU33Fv1
SHvkuAH+p8Zuq7E+1LCUY0PjpsIbbM9NWLKrizjm5Oj+M8iHIen9ocoJvxhU5kZUaKu5p/WCrCKy
e6zX0E4IEhR/A2elLrQXro/ujMDopyxBD+zH/7ZLTzVJYTeSUhIqv6mpDWIvZHE8elLvufdXPV0L
Tzb1SOCg28SIV8pkSi32aYxgq1Hxu5n/HUpSH15PLsnW4GZZol45LM6/TKe+Cx+W8Ss+7MqVMTg2
wVwwirVsiyjOnuZnxdNLBw5ZMim7MiEdyzo5QC2hWm+tG3W7cQCxKKyLH+p/1DLizAQZOxcHW+11
rWKW6stdaYpVGnO8j3b/rHt5SkyU3OmUoll5Vwp4r/jTpsrhem6rHl8TEnA2bvCsY+M7aTvxSBn3
Ed1ImvlHjDGN72pGFHxw66s7T9ixkzHnMnsVC8m0WPRV2B2bku1PbyMf9lqJvx77nZ7AxTe5yztH
wtLbMTpZPr94mEqDV82TgQxrfo0B0Lj7wcfHjBNJT7aoMO770blaLuAg1FJdDdzKZ1DeL4zUNZY5
vr35e32xekbij5rYQCA3YIY+zdHVcCiHIWa38jGw+7vv8MHRJoT9ZmSgNDMQxIWZUJSRbTcVYTCQ
L7FptEDyopAeDA9WS3+WqrtaRZtVq/3wL3QDNuFrRKs7d8JtdR7o/A48H7MDxAWFryNVL8iXevFG
QoKxc0emEGv+UUZSIZ2mKTLDbRQJi4qyfz+A3XV40kXVZPAtRl7DpMSH4EO35nST3av/FczGAajI
MhRw8vpYVWG7xLTd5jnYGAqE7cCzB2m4L591S/8jlGlSDEccHMCQ1oSnBM0wyck9KeL1qZiOlr+C
QEizfVWGIKzclc4Bom4mvkpq5CqB2trOPkWqv35lMOMykigCVqsMikvTSd7iFzocseJbq724iMFk
MmMFUDBrVe760KIJxTMzJfVJvs+0xRq5FVgbrgZlRJFXRHykamKkapUUWNk8t6NnLqF9X3rPShcr
72bUwjB/ObAYwtvyDCYta/cgyh3QWC13J+DdJ/D/Sn5YS5o45mXVfGB3iIGfvyJaBKhQrIljO2RR
mYYSzSlPikdY0XdDqASkSXhGxf+su4EmUrH7ClZQ0LBy5ZVYx2vbWm2F1Gt6gY43SDQVlBPuLXsh
I/fHVPO7GGTP97QjaqbJBSgMoh79LCLQtvbTSNb93M9Pmphq7yEDhlmMg5I67RZAkUvXa9LWbJHB
LJrkgLRH9gZWDgfhW0XQijqsIaDI74xS503xmsp+x3pjDZ0xuEm6MArLXbql0T21fqOwLfaagKaP
4npzZ51XPDDKaRDyyG0ew6CvlaI4WgXI9+VrS6nwP0RgGv72lzcJQ3UOHfNfK1AUlPhBEMjKeU30
v4Jp3z9uY5vU4gLJrbVHRLSdY4Fvm+ejtaXP3B3N9gzZ+4Fo+t7RJfUZLE4TdeqlSGn2unEQSLtF
P8y7HGCOyPrgxv9ROmNcRC6h1hQvCwc4KgdXkV91UWatqOH2wdzcs4VQyajeV8SfNFy2tOcMVxgb
6C3KDyuaCrha+nHdma2HvcEpKgzFylmBbPqUhWqowqlmPLtdO72PPtOpP89ED8CnC3jEa+PRgqNH
ALbqFS+eFDyQg4sxck9gOmMqrgR79QZKeU57y0tuDNYCHssLbYiB8G6v7IfrO2JFLt6Bw1p/xNIZ
lMKhQHok9D3ZqfqW0aXGmskSL2WQ1bDRD2V07r0UiypIgK0B6J6nrHNQLVgJoR7SFUNM+Huacbfd
oLHOMwLy2NSFFkO5jzgG4uAyJXPr5M3t5ZLXNqe3scAy2BmQS5lguCxCsr+RA2/V2ibrZWJzrVGg
qraPBHVrzhAyeJH2Wk8TDS6doGjMpGAcuPWUkO9sKziwvBt8GPh9ZWD7cHGFsnKN/MPQuaBpk1/c
P3oTZJPx2ufguQUDTqrFUj3Tq+mdwXv78J3mpM0oUi66WRikBf6AS9bZ2XAWn1eIFQQFhvtLMebK
lG2/qVxr0FHIXZ7l1tYbaMpKDhIl/fvaa0P6IlO+VTOwrWmt/CnRkwJgtEW/r/RstBJsZLvtZdgP
/ckTjO4TE/LW+AQGEFvuxjdehiI6K+oKt1lKnMvKwlHw8VY+Dzrkz9JJgZxNll1Ea2L0Dn2+QiYk
MlDb9rIl/mvkLaD1lLy1VDTKSnu4RxM7isdxqsV/nWC5ZLs73BNSuG364denu+gsr9v8IHxVHunL
zE5YC+xi9FLQubV1DAk2L+g2dg4MAA61EqpN66Sfp3YuxYeizdK8lJN18fklJjHlHlILTv5a7x7y
1OX6w2zlqGQFZSXzchB6WMeGSXnvPRozQekKimV78s6EYeRGRccTpSTSrNVozMGEd7FKBRpAjcs8
YQMaCif/8ATk1R7Uve6p83sfciwGLtD91zrnaXyTofmkqnptMGxh8pDERBp0wAOdAAqHzGxjrXnx
H4pO2FCed26u8cncnhDFb0TUhH0PMS0nZ7CbEeLZowu+NdSZt0alowRCyw0JqSMfY9oGVq+dt/lc
eRHBBPtUHljLwJIwtSYJV4lM0f7qWmndh8n9JXgQyZBalSZ66WdqYw9XzGVtw1SU3UO1jRVYrLls
ljJIGw8Gu1XDtom17Rf7dcxnj+OYUB9BPXN34LEEH2/RXVNiFFiVoo96kFh90e+mhWO8USvXAjYQ
cqXfkMwupG9zFG6xbMk5LUmVleIUkWFnZqNfzy/3mXlvMgAd+ot222GwSBBQm4u0wR3ekQeyfNzb
P1vr1KjPYC3DZaFPFDJb16Q+8fUvK3r9MsB88c6nvuNqis1B6KnNhP2QMo+RCIPf+osyOz5dONEZ
/MbImk7PvnyIWJZ4fK0KjBeaAfX1J3Y3lVSLEL76XDXYHO2my6o8LSB7bglRYRshkbhStan3cobC
tqfkTvxvizFgsZALWoYJTRhllOqhC2TYmr0pcOhGIDTAcJJO1Q4CcTzqnlGPC/Hm8wlt7Xl1o4Yj
17m/qi5kpnZ8xLu2pnqaF+mhR3yMK6qMj+ShM2N/zT48BaQPC1N23kihKOBu6LeLjpOnBjKKmrTI
n+qTe2n/KLJWW/RygDAftRitFjnuJvD9pCfm1wTKwe/GsO738fZ2+YgF8SRfaeSoSB6hE7ZgFAZR
Nqdzh1iOIAMGoTocdkWjDq16Z9vo5faNX2aYKYaLKa/AkIwkW5jjkV1lrJqc+/UrSvITu+TJIa1u
lM+dhwuQYEzXPAIVM2M3V40rNTLG7VvlobI9pSRYyTOyNH1h/osJyJ6AWW/74vmXdGLttMnd9CiP
lWioEMjVKpQS7RropEqlsKNrvCa3PRgtY4ejO+vjKEtoTE3mhOakQkFG8q/87AL6+PLhrc91B+uZ
Vt2tSUWUDH4HVDbAuT/XyvFc4UMrwZ7dZsLio2LRXID88LObOAZn4ieiqTErWafjg8WgjeTrbws/
wGoggqYYX5JlPyybqT4L93eqWp9omLjdDG48FJeBBH6+ZPbRVRf+v+b5hrSSfzgv/Le5RG0eEuBy
iDQRQxyShCIAT6d6EJQC63Pldft2/jJDD/tPTakkb/HH3K4M5el9TiRmQXCrzy4LKR/VZbvqDXy8
vPHnWoIpY0QU+9vbTny/Kmc8iR+A5z10U+huQgZHVnaWAs9g1BYIJsU+8ba836VwvWs14OQEGX4z
COLaHvWMJ4SQNGPI8+JcqdnAOPVFnL4zqhWVjyT4heT0qUEubtfRDUIMeLNpNt1LM55GIIXJpBm1
q/APyZX4S6oYP+o+aIc2ywLrEA9pQbrmL8VUjBTHa839PODjkaqsNfmrFhOnIPJJzXV8jpSwEN7/
TeLFeId+yr56HQtXMFutBYsc/ND76oy2NNOa7FP5daYVCY0mGhR2tBtR7NC8YeU6V28qoQLs+2pu
PQmT/XHyfb768QGszj+QFly4Qcv7o3NjK7jC3Ad4nLOPOg6SFLdTFDnESJWv257Sun5UW51Jp37y
WZF0h41wtvMxWk8A8VhM/f9IdD4TpqMkeXqwURBxewbSFs2QGmsZRIMtMaTbVoK3Ok4WxGu1DFtQ
u/U2hsKFEBfl3/iyXGZhkp9OIIgp495UTVNNF2y7TmgF7PPgt8G9LuDZg6+bG8HZVVamQ0G2mhvn
IfWSgu3nDwrdUphcGjw9fdQd6X9rK9EsQ/ToAvpsudxJg6mectDqkDa3aRvUBLMK6zXtYHyE/Nd1
h58+7yGBmi4liWQ1NAuNFoDwCsPqMFaqUmYMjgz8fRZw2/Lx1Z350J5d5Qpcrj+ZkmY95d2YrGCF
dNxGyQnZCSRs1lrDeqxOnfIkesT/gE66S8TowedXwjTizB5G99DeFJL9Ar5GykRQXT6idPMR4iwW
qzijP81RS+UTG6Z72gYLlMzwATdPMNG9V3r/QttMR0fd5CYrqwJ3Rm/JzleL8Qdv6wFTLjYIwkjm
qVQ/EkU4K+18RH673cc5iIWjDX31XmnLoTBe6mC3JqD/wqBwGweQ0MVxieUOyZD7tTMAXJtOUnEZ
iU4Pva8E79wtEQVqu3cfIixY9lUxD1fnDUZwovYN5pOmVg35INuifHJedzZg3fMUoYwbzzkz2KEt
ZdG0J4NmHKbRh+6F7+AiX16fXZbpYE3l+rIN0zHAERgPmDkzgTG08iezijYgTDEkNM7iK7+8RObO
wJFG8gQEo5eSp2HaSNQEKdCFCRWE7YDFZEjNlpUc5w2wcwipyo0SMmWH6dihVtot5pH8xMtPhCeA
fiedELfeFhwxECPGFmqGK+Sh2OoEJKDdlZmIJ5oP/fv+eiA9ZTD7WjtyDbVRpyAYqE9Yoc40lQZj
kGsX7nXcqw0DiTQyWOm0co6oKyidh3ipjtGiFz1aSc74GmR5idzD6stGdxXkuJDJ+6eY8tkqnBcs
PetgwX0SmBKB/u7wIZRPYOEcqWu+OJx6UU7YaE8HxvcMRgGElyUG5u5Fw4H/qptUbimDutEDs6c5
ARnVEMFYwXYHUBzod3X3txobjHUFmUZtW1PFB0+zJw6Z/PtJYEZUs0nVm/i2aUP+qbc62cB2vHbG
x4mAwiDgSIA6oiTkl+ekmVA9KL83k4UHqSeGtT4tOrlrLcmPVuXKCpvGeMt4Vl4WR6l76dKcTb+K
e7ehNUJJsiqyOUiSr2s7GYPsas7lRpaHa4wBlpg++QTI7CDXmXSWAdO6nysg/kNXaeldJJ0bsSO3
aIfBfkO3zqAZkqVxPSfkX/8lYTXLcJ6sYnljbAFSHVXpvkyTqInOEaAMX2eJ05JWWdGCcu+bugk8
GfKtkMUz5aaZi80GpXCSULIite4j1BK5pmhxMWSKnOuc9pg7QS2S/AqjzABrVGrl1h4omLyjE55/
F55l2sFolhV0Q4Hl+C/I9AC8LcAYnhOObrszCZFDreRA6Z7j5eS93nXP1s2PhJYHFXXI89ObtWtH
AVkM1RE59+zWDlf8cT/TtBPTH0PKvdvdINHoLaWTVi9uSiJcbTYCIJi0oezpjfVHro8yopKGtcBT
WnZqw/tM+2MwNpIIjLPO6/xJtDQWKTEHhgBZWIQfBrkIC8X3HZJe9TxyDdiveOIhDXv1TeIzYliv
PxWFgxY5gg2OJQh4PL7HniDKfPJcEMXS01P7DyLpHTqgOXTJ7ipyvm4tVvP71rQMqpiWfAobqRmY
L/3xX4AVUMWVW9Lxgk5TYHWbhqPRwRtvQIuiIYe3AG6aL2i30qC94CGwVMm2akKr8Ary9cRDHbV/
J9kHish2ve4YkT/c10xGnPL5zTcPgZZBQk7yfRK0KIF3ehl/sg7WGrFYMqCpFj3UPW3B5jHV5/bH
HdPZNmrU56gMjFH5kiM9B6RxY5RsBfsfEVkICLVioXTTJr+7lyNJjVOyQ6+y3+AWXPP+0cbGNx2c
PlqJQTcp7m6i88rWHTAw1dKbIcNmN6QaDgAx13Y7r3rzQyCImIEVKMAwiGd54DJU5e4uBGB3Epsz
44+sLt9+gwyayY4NVkk57JV4URu4GWz5dFRzxl+s6nBfy6ypo1XnIbjqgGVqgg1n2FHxiWNNFNRs
ks5EHJnAv1+zRRv1FxmhRAucUPacDE10woZPmPl079R0scWYd3DbqUJZzwK0ewWl3nnkHEAo/l58
ukF5pWXGpugsGj3qTBuWf2CWyK6nFPl9P/x0EFoDgjqxscxpEczuKZE5T8T+nA+P4Kea9V5vwDV6
6zaU+x44zwNGtDzu5uSv0PqvPhflNFjdnBSM2rc9tnxwDRu3fXkFvwvbv1byXdDeBwFqJ1oxVASK
RAfpeQQ5h+YOkuIxpjxnzhvin1BmaFyKmqf9RDfIE9Bs8f7jYJG16yKIcWLSJMwd2NngIRGdn77t
Q1TUF5cGHKRyHfk+P8No5zqhP54Ve3IvRn5h/kFjRrkLF1W056As1LURAiTgLPrwf+x+WFJiarLI
94JAZz9fZQn2y2T6mFuxerkbkGsaV/jCR85XVNX5DEx5eyDroC1ThvRTBdCs7ZK4GpQ+t/aeTaRV
UlztC8KNG10li116fpqhi41tTDrrfJ28otfy3h7Ve3HH1f9ZgClhV0oxbFADBa5M1OnQhjNYx1Er
qhPh2IR2tSPb+RlycsuioCBs4wdL5Ramn3rGFS0mQ1dhDy7+CvtZr6bDQ44csU3S2ryEC5eF8sqd
XqOIERvG43Bj0ewXn70UgiNenVwSVxiVxBmdf5t4feMPaO/0usZcWZ0j6h5h7UxB84mVKSboV+A9
hiehxdPbB1MHDdLsHkLcijPXXbwAyuK8vSYyJ1wt+4oxyee/C2vSQToWpWsuIb6gGbi/hMmlRSEg
YsG0bkcJBaH+ZrizLbR0cXOijPcN7Cqwss1tGxhjcCCMIRDc6qa3NFgZxgx/WQKfHBJFL4lsmvSl
AMbi2U+1B/MGlBb+ljPQrpIvmccxfSaMEE1AcYrKZq/rAhBqHB0WC9AP2sYyoNAdShzOb5afFHSY
XVa9E1NVG3N8sJKp236fdV3I2ZVglm5YnK3koegjb09qYm3WxCvrAlRPylVJWyfEDQwf+L1BK/cx
t7+tT5kAiVd7Si4Nynk0rMFxo3nLjL9sWe1vw8wx1Xgycn3XuOCaUi1umWSPVuqd6alarS+MqiZx
dM/uTAKIaoK51FgXVaoCLtfyrXyt7Kig6sY3pvV8dqYDmkrLE9hnP9c6/vsn2q8l42XRXEgh57zv
UA83UmvASw2V/pChqKJZxJaaBm+xoudQmbtiytmMfehKgoca/f7GVEo4/NGfuqNMXT2WpGOht1BU
Yam8e/Q5/2o/u8eh+4Q0J5EUgHQsks4gzdw0AI1NtN2F5V4pMhziu0b/sIEtMJ8Rz+KC/q0Jm2OA
bv+vMJb50t9LUeai8jjjtdfk/qtalI5cBIQitr69Fv26OC2FhYKFiMVMxoz/aYSy8mW8TiSoLugB
Nohzu/2nn8aNWwUPsQ8DWY5LJfK10BFAxTQ7GETLth8q99IM245fti+iCJvjC3cop+sVSQPY9Vwp
5dxu4arLeyQ8agaSXPFHY0OQQUW4wp+OCwyZyH9DpK/PwsIZQ96jsCm/EpDbCpVw3plVMiQ5lPmI
Spis5Y8sKkLlY079exJ400JwCf2mOJXpBx7DMpp6esTAOD9I0aOH2KNk63Rgg9RfnZtEC+hB1N/I
Y7MHZZHf3YvwQ16M2hCrz2+wlyfel2dEfObJ2+ssKVgPd9rm1qNV3ym8cKSzV2CH3OU91p3ZCY3F
quYklAOGDdk8UkJd5YPHtcbE6xKHBckWG5KIJjlp+4aM/dT9viArsfJnWQRyX+yzUh3nW6UHPDnd
bnE6WnbYRbIcmr/d2ZCyVkKXITWO3yJpJnOPcx2iryXQHfo/OOg4GUL9dh6BJcQqH+w2ZuszdEl9
BrFw5DKgVmZW5CURD9YiKFFwG7Jh5UaIn/D9BzDvMjknMlPv8mLmqn2cK4MhbOaXigt4jRpaulFW
rOmOoJqpluT1jOOp3W2ltThK3pTcVNvVJxEXJUEfbmLDO6nyCOrYkJ96libc7AnF0AYQ08ok5MLU
t/PAbyY2tRmGSHfxZvzM2pqmKrlFwi9B9Ioa2vQGumU0T/rQ4ob+wsR+T02R5iYP4aLeQ67vQiQ5
JC3x1kVRTePctQL4Exkzmw9DlVPjLT3C/Y7+GFNb/FqhvMiUuYCeu1LL4NwTvYPdj8FvNx79aix9
uv2CZnBJw+vO+7V4SmSgHyGVEOwZGR+8FrYI6nTA1pts/He1tSV29dnqGf4hoqxkfpr74irsprgT
sTUgwL9BqHn5d3Ic0y2rECZeee2hUjejd9PCr35Vh3AQ5r4WWIBx3mlX0rjJ9X7s6Ou90jnpEe9Q
ylSwSi3XAL8BS+JqC1JhlSqoM1tBoBXDyq3ryr/npp6GmjlCLP4mIoNqM4AG/fkQvRI8z6rZe4mG
pMWD32Se9lki5b/vWvqc1rRbf6nUXTugfVy5kfdTediG4dwm3V3vZhaf3EF6esfp3iRkNcOLxVSG
G82SGIYZDl0RuZap27xdufNKWaVpuphkYY8v5cUPTOG5LU+gw5tgwRY0npVzfaFDoC6fbJiWMAzn
JvNxyqOXJ7XCHTlaMwZnEF2LAAWuL5D8PddiPzaqWU6hDgkbl9jPs3KECM8tg16kgmXiTmumScHr
9Xa9i510lG7YstcPjjOp8jwcJwxgQUZbFJ0k3fUuk3qckEtnX4nUfsmP+dm7k1rr2gbLv2WzJBny
h0Cdd6ciwWBtHqReQtreYi+R6IVLUWvQLPSVteDZqj0LYYR+xt9gembFOW8CYJqeTT4HracSqQ9Q
8j+2A45pEn+rx0RPOg8Q/M1ZALMMlvrqe955hPdP8sVyFe9mZ/vNntTk5V6ujBgrwp9A3xc19pCM
ndmelZnZuLQG8Y5xzfGMjQs8TzcNF+BzEYDFtH/VcyuA+jDNULqkTuSYg9dV49mklOTkQhg7qwt1
WY65Gq0eh0DlUxQEZrGIDaeJCgUdOhvr488FgGkPTyVzz4RnqQNwvUtdFD+Wea7CE8ybjD/m3SNC
9d7WZgG5QJ8PyvzW9hEK4eW5BeYGL6/0xGmVfhyBZfzEptcboc7Qd33KEgdFp3bxGqQGJVExt6qg
6BzRA6SkN6WshKkpOW2rrqYPNrdB+gulK0JK5b/kKuerIdYQebi4TrCjo4zP7OMGv5Q1R7NN5O/4
TFdmzkR0N4tnbi1smmzVt512yybo7239o1iA5xdK9E8HHYRwlE8avp1oDKcamG2y55v9XmHUS4oA
GI8sJdGJV2G+irizytnfBoFllAXgRa3OqjmAJi6irHKlawUEg5vjIIekT15+L176GkWeyH3YvOC1
WjXOMeP211KNyt1P1+Cr8+/wwocpyCZuLyY3FeYKcSqpBJf/na3TDHBXkIlYBGSpidrqEaotUNlg
IkvacDnncpMVeZfWvjG+4xT9Dm+rji7V4eSFCUre9W/6O7C/aaIot1/p3oY+wL4l8s3WBSJlooDw
2rl2YVkg7Yuuk+MHduQ+APTnW48NXj+QvYRdYdP1qOdGl2muUd3lSVlstDCoLt9Qm5JQVHElkf2O
C0U/SdRVuuN3lgNbUE/EawfJV6lITzSAUSviMof2x+aEsYAod3G/Vkz+xRwDbDHovzzafASi4ddk
BBxfSc+SzxnM2SqGmxPkxq1sTRP+4HLBToFiTtwZHrEVSnpf8/KBDEaFapU+21yQjann12f5bJPL
hdvxzUNsMEVN9+7MqiWHa8aNzXGLDvLmbaHdp0RKjq/HEvJiSle4jBVhU/zQm6EFl8HhPd7kOynn
HSKbaKoQypIVwyeC9UNks8iUuz3RjQNX2kt0aVCESpERDKkHV32BHg2epcK6+F7znCqjawFMrQx8
tT9kETfrkNkLTZXT9JI5KpSL3snQGlezMRGdHjxnBrxBHJxVA5ybLnNd9sk6uQkjVKTidKX72Wa2
IzNhJ8kLo7zvmtwuf0Z0owf3N+fADDT8yV/nhSMR9+SPR5oPtHlnjTR/neoOCSd1uSh/SV6mh151
Q271NKd9G6ff3ntAsqDCLuc8gTPPgpeRGijHJzOx7Mgiquweph3zR+6ycaBjOqnq8VBZteiud9a2
wPFuF7x/pQmyQEx218opkEJ4auiKcNKHuGanmSJsjoYi/WdqKSCKzJV51f0bRGkaRlM9l9NsHsvo
fE9d9T/X2y8aSS2+lv9H8U/TG6hIyIQVjn3w2fgnCtU0dhMo8CG6XH3YQKtD3NJjSvHXLXgTLL4i
KyAdSbdwMZE1PYIJi8y2oT3Zc6Wqxj4+pICKq0OobrFPBSBRv7UY8joHeV4ItCTZBi82ebg5CaK0
SpA5J/KK3Ex8aZZwy5r/c6OldPuuUk7YoYId4D7s9lAAHhkfGmZLXfecQM/nrRhbBHRsow8wpt74
JyPxpjHHAXO251QO1ryi08v2+mSd7xqwVaz9gF1yppKRMTnn4Odud/ZtoKPQDQJ0Gaw/+aYPk3JM
9acAhXy2uk9rK/tELZJh9/7SNSlTa52Qwic+e0NBfISSzzmylvl3G5di37uUNIIRtAuHe2avOHwv
NAS3V/BIlL6yBU+cPrXMlAci1MrbrXZwrwBSCnlSjAqubK1dmmNrocyIoWRhjAOkbey1S5kiWdB3
lacRIh9ovusLry/CNk0aql9zbCms2SJceRdV0YStwrtgSr3D+1DKRkBB5lb9Dw96A2oscKSWFqba
e6+MuDwRYrhlsN6W2HmGxF57ftNRClVrqczDtjZGp7KhyVekstrKdqpZrTNS1nz8y39CAvhPXm2Z
akTeKO8TVjyf+y2Xcga6kbqCG5Eyalfw8T8Q7/U047761i4WEtSbOuDYUNhBYKd4Fg9ZGUV+uFaS
1EtyN1DLZG2Jit9TVUbof+EGscpEDQ5QqQFyk5Vt7XORi4K1srGUZZLpndT064IobBLxIBwprT3b
6RtqZ8HglBgD+ko/DltYDb8q6S2uyIOsBULeSEOCV+aeXoqGK4Qys3mFpwtIUf5ou/OkbZRckGT3
L+7bCps+WYbYBhLwzfL+PR6ekI5iiBkJF+RLU85oaC8blu4y8MSMHpz64N80AQRFQSBT21U4v+FN
oJEGAZSidyfGuFUw85/J2E+iXqRo96y4Vky5gGei0FjqeBsmhC5yYaiA/CVLnQNXunHlxiM37MHk
R3hFX9S2Mhrfpjz9L6Z86iMnYTxEjrmwKca02wbt3tknusphkg6foohoK8RxhDLhrXyUdHZ5Gp9C
BQKkqQSAlfQOJnDBT+XS0OGNL2cFrHyy683JFxH+vwudzk9b8VPcE6uO811IdTTdTcDgRsN/Xu1N
dP2tpe2tKbcLMTGzIDVVhpDaNE3Ivxbw/UuVBOUNCfxHPik32T32pZq+t/GzdRw/VZtzYLvoxSpv
7BgUdlhwmF2RnGEj5StauyFFi8GtJWEqXM3VG+9VaWvU2zZ668ooyxZl/sDWu/fPR9qxbuo4PM2n
XedSF2gBSA3IdWozbtJtjdibts7dI9hBsNNbDoLUOwNZIZ+sXfsccz/0bt5/UaiZ89nsuMw7M366
Bb4eCoJXDcrBBaOU98tVvdzns6XQ5tfA8883mOMHWQJM/nyfaYpasgkrGGcKbcnSNJSgDKO/jqqz
0Y11nsM1Bz/1hjeQYnHxuhH6PHiS0Go0riKyqjWfU6xXjQRU7+B1Uo5MMlhwtkx4Za3UAG8Zj9Kh
xcCz6U6VEhKKsb79g09mi/45mf4LZ0h9ZK5icn0hRAtZ9n6xClFpn8GZ6euEjVoEZwvHP5znqjVd
FpdvYt6z2D2e3gERQPqg0yaaSHiXWSpBpVbp0ye8KkUf9c9rWFMcsLhCGhzQ42YjE3zv58/KuPzt
GRrwDw0eFsejqBn4s4TBrNq1RYSwGizpMhQpT+BPvtY4erI74HaOvw8cIYENCDhR/iM1u2O76t3m
03/7ekRdKnzOFxLfzlGZDbcliHDzm8+paUnCFW8gdOipD4igUC91c7SyHF/bFc52LHI/THMY49Uq
+4QA7A4tHb0Oqr/0WMO5SwpEotv+OStgEfljgQ3t7vL+xKWC9bQdPA2DU16azHkiuYdUCZ0dEP8X
S4EeVCj23IWp4iQ7oM+ebN8DDeNCADObX0TQur6o1qaTjbaa5669BX6fpK0bhO0qsWZ93AaeYs0P
SA4Ru2SiP5NFOO7jEp4WfbQ88CX59xWu9WvBJ1IJt5l99doK6z+lt3VpIHWM9wXsyEnkfZmy+eR6
2tCY8yBfVxUXSCO9oIIkdY3WjD1nD60/NMUZrpqdUm4anrgiLg3PgZeYeUE0Hi8013Du8RFGzzVC
8vElxvsIDkEh+PtDbgtixiJnKznmr2sQ+euX8B3tKGx75xMG3hZmZHp+6toq3cLLTkOfzO2KD0pM
G7Idf30PBA2FGKtuZ3uDlreQhFsJw3Mtzzd2u8SLlHz8tnO1D+ky1D0AusMG68DlVzsDXz13aPt/
+bMdlWeZoKQEypu+I9GS008rG9KPb6EPksE30W8Im71eUi05eEgjxskVa9uWrlXuHgcNHhF1C8db
ZkRLT1eOvDH40Gv/TbUAs6IODNBTzFiORZbi5YyIKlsrfTVyRdPZ3d11LFCqsxCdEDUOfTk6T5jG
z7kaKA+WMaE3/UsZw4UCe7263IAOp4k3lIoQ4pSlFby7X6OVfLAhUYNWf07w6y/tr6JvCHMQscyi
9ggIyXemPYRmf1hEkgR+FFfAEpxmZLhhbd+/VonKInkyZV6Hq+4kzYrmac5VmrqdTPmgl8cqkJVm
8zOwWJh8+jAmvBDmFb8rUQ8Cm3TX3RWzleJtZ/kFQ0GjoRmHGjLOMuxEe3oRBfPGmH0abOUfIx2u
e+12wqiDI2cdLhiMd4ts8LoTi8BPq120a9Nuo5jzJ6FAErd2tlCOsPPssyagnbCFH6SUFpj2gRNI
93hqmnz+wbMxH0Patz6oxa//V8kBZ/9jFatYukmqPg8GJs2VQWRYi5BF4AGWJ8Ae30MqAvncmcPr
cNOrBJZ2kfBHn3so58oKOSKFVJKnoZPxwgFyIaEnNjLuk72eZZTAFES68D0OoJOS3UgYO+JlAIpK
e+n8DB2656rLG6b1uxWBVLG3vzst1W9/auiI9PealKokUTHOxtSRqTY7OIpPRLMm79SvhIJkDqeR
1WUHZu6klmKouwhJWvgQC50+Grfv3iaSxTJ+kVaR1Jv7Gn8yEmlNKH8ZgNVRtw25sHyWLJDKpo5e
mge2iWQjvmWQ41sacahY/SoVZyNDyl9qxHcWnnXVqN1WxA70RIMjQ7coHXZfwmpV+eaIpXIBvqF3
wmrKrA/tvDpcOIeQvRHkTXcKQezW8smLa+wWAmTJ49UxwacR+M4F6zChYfC8IdXmxApm3dm9uWqX
2s0wuGQIgsNYe32fGFA09PQ+aiWCEdH6eOa91PqBg0Hdz9C6XonpOBRpepu6wp81Owda8msdmLJw
76QqRTU2MYfupSa04vxvGAkQkFMNTrzMDR8qIy2SNiNSP+qSYeLYLhGlZZ7peFyoP+Uy4tUCGy1F
Jknvn2ZkcBDuNyoc3xDRTSAkOWKT6LOQqrhqjTBFe6vR6mA+JsBajXZC5W8noeSEVjeG/ynbCmOy
bCDzMkHe8QValwhmSjxgPeglQPstJfUaRAceMrI6LUqaeXvDA4jGIBZW0zfc76O32jJE1qVAKoOk
sLzQYZy2wQhmKK+k1Azc3NoLIvHAmnYsJYZBNa2/TxeSChw/sgtOCiLDO4YTcfPjMaHpTjf/Q2KM
3/Ait7TXuiMPoNIYINwVLPn29OQJGL3J89MvU8R3dFNAFcvj3hIEjeI4M4WmMbK3gUIGy2NqLreJ
NS1paICkOwOqVCiQozwHGlQQ6vA9MoRhQuxo3vC7niRBV1JmmmD1Us9XQbgl9UPO35jmFyPiYUFy
IvnhBTc1cI+MhV4FjE9GmCE5mtGW7njYQOzAxJkgjeagNMwjpmFKoXel+xRY4Bpnx2KaVedGZCXg
qTZPwwcWcJXMF/2AcKuJuo+FBsZ+jTEw/Am0sZ4KX9Rt2pG9ILaVbLdZWiXcIu9xbnl1+Ld4de+9
B5P38IzqPFoAZSbq/3j0+HzCfctiA3RSOuXnPZDp2vNLaoGUCFiwild98fq+iAwxHD+khAFMe/6B
SI1lRkBV3LAi5ymnuVjTdjowUx+Dcst8/Hx/ic124fCciFz5QKCkPp9YR0WT6dFVeCz49kWtUEKY
3AmYvOl9d9yB7kxRxT/AC7BatDtqZ0hQ2enaI5takgNJUMKoFh21DL4N8QKROaOS19GLbTk6SxbV
QplBF/yeKpfJYcxcnGJBRNV97ipgbVQA1CNlAnEFCG/DbgPXZ39BNSfUKEoZM4Mzs+Kg5a5ACsZa
s111mv72Hk0pWfmIVMjCFuFpO55Kpy54W5w5TjblyoSxcLv2eRYf7lKsZq9c9pl86xyFqZZw5MtN
om7ooWTHfVwqDozI33bCQsysTY2RR00XHyTkLVA9Mi4/lW11y2OF18dYV+rmuUKjHukQ695H58Cw
IBM11WPxN5oiQWWXAo/Xve3BGzPrPBoc38HRA1PQLtae0ngkkddB5n7AIr/aoj7bxdJ6pilpqgxb
aBB7Th+QX+yKNgZ1I38g+14LAfopR2i70JHbDA8Mpe7x6rSsV4i92dluGKP1wXts1IxBpe827n6L
Pu1l2SHuRhcOGOSLflhnyAVbHQr6UczWfqe6f3eX/PwFGJnjjM922DEOb8oQOu7VYt2ol7w2UqMY
PXLAwnLDhe5ofQ88QphzzTec8xqrv4yuLybKaMeyD8Nrwd5Fb5J7W3WYCktqmy3awFrQgtGvWOJ7
uXjI9JGbstbX4PYRkcF4JPcQd3J1CJpRLZem+zrbEhBEYtn1FFIzFotP8tcvUd7oullSnQ67L+IG
nX6IuDakJGtACjPJq7aMqQps1LoUFegTLpotq/h/OADaHUOOar9F87x8+AxqZdGQ92VYrw4hWlBX
y9nBMhyYzaY4gHAEK3Jvq+qDTdhuuGGZGfy0AxkssyIDG4dfKIosWgLbQdlqVYGCBaVQcJxqO+4t
5d3v0TwNPAM3w5NAsdD8weHaOM9dwNbEePfE7SPfrGx5sLCDyZRHskXvurobhhQSNKv/zbwsc1DK
nEjdjbNgVX0aEjDhWrhcF3bjjZuC7SEJfPlU91QmcWdLkneEWM/omI3A3J3Rome4ZzWDkyyAazEd
3gfsMc3dh7yIZirV6l1NUKpXOennNdIpd8CUilFh9bwMODxc+SqHghg0uo24/dGYJoVo8uHPPZ2S
5sr7tOg1BL/xJvK8t9+izTFD5uK7KN8ob5Ap9wez2tA9IpJ5ESGuL1Dsf4+3QoCdpALFf2ywTUys
nTa18c4cPbiYMrEISsmD+qOPH570sUhkfAqlxB6MWr0uFHX2Fh4tC78LjsH596TUx4uEFSH6O9uY
LhWYb2Z/z32JPYuLkWJIPLKVZV6kyI3HUVpc0+ihJ64uDEpgytbZIRzm9suviA9LF8CUi1ofIXY8
dqbcm/BYsdYCKtHLJMJ11M1e8aUcP5sr4utwirzNO2sWgBJglSliTidvg/N7AMT3/hQNv+KxEeFJ
wYekL/JtR5DG9VSFVVMkJJaU1EG2ukz93LJHrqgZrF6bxHlnIB/d3554tTC0mVqAurS2yYn+1q8/
I9x47vQAhZLL3DiFTYpnnzRZ+9276OqTZIGDKoWPC4ZWL0/VBg3RznUfG5MzR/rpRozNK2jcn1ED
w+wy4fxlKk5X2YuKD7HLaEf+CeSUUEvlAXO13mqkCmc6Xim8Ahw9n+9+3Tf7YIPV+PiCx/F5ukHj
vGVNZdrlbSrYFaLln8A6M9PLSzCC45qfnknMVq02L43r7D7iJmiBsJCm26vA3YJP/Kn2EOwYvnik
AJeTafuRjTwHMT9IAFwx2HeEG4vY69EzO7hE7bsntWGrUJ1uISLrJVYaFxErzqC+Y5GQpA5FrC9r
qy8919Fvego5t6HipTwP8HkBM9aUZ+a9QoyF4Nae5wr3/2OEflDhlGWW2BmOJeZt1f9UsPMZbT6+
bdUH0nyqitst/jfM5Kc6Vbd+npLIOGq3iv1Vas8a42UAG5iRdi3RjDKBHGOov7MsCkiR0FNWiCeJ
7VZ3nC7sxw6kb9LOhbEpsWaXatX/QK5fMigfCZ3T8Y8D7GewOjGw0ray9oKfd96GsMaH/6NdGYHM
KRLbHiAxbsWbPCNhY6T71Mywe/d1lxSMYAI4mHKNy3zIWdGEVL3/O3duUZmFqkZutRAoCR+w+wgT
+Adpao4dkRnr/cIgIkukZQcyRcs4eU66G3gQYanJWtp/AxH5Zb05eew/MDKsdvInfWnIeaRwSOnR
cufhKQ2TLBkKx/jXurahfhkSBRGnfgQ2vETzBjX0CJaz9m892BCtlzLBrcVkYrNYaIvfTSifCnkL
IF8SLfcXnlHlucVWWBdJKeX5O2aA/FmbV9or7zyehcesgqrG/SpDWN9qTdUyXhdAYtIG2/LZkYuO
piXCdqsB75efgX9LwbduhDsMKv3/T4VFxdffQqCZJv9ZYf94GfMC/8MPqZ6shq7if1LjrcGIrngX
IYNG55ldyU5lYyd696RdKWsVlPF2b8sFZvDr7Xn26ekEawLuRIIdiKJEk8VqLSorssOCQquuy4gJ
lyEph8xjXpEomqyihhSg/629sFcvyFxor+hiLHOWIHB6F0AC4AB24j2qdWeQ+1ABmXEALNn2RZiV
T7+Fo+j59VBN3bP2CIp1GNL3PAJgRvRioyYT9sTz6NyfFF8veMNbfhURXc3JP5XcMFicjd2QrpKL
e2vYr+wnXRI2XFQyOMGDquc5B4lOHc1VnFaXd0YQ9XngtBPZznYZq28wL3kZzVUAjJlLwfL/oIjL
trsG1QUTHADAqfYAtMsk+HlGbHyz/hpkDDYaIrz3XblfAPqmZl97tA8sojWJRH6nk0ElXmzz/mCX
NTaUe6/JMJUGM860+KqNSFTZfSOnVo1JgMsN6icqUzZowZDZF0MRTEJIeOdT/GmOrdnuWcg9T0E7
9y7ADbm8ixaa+NtrYLq0KcZZTNcFl6z5E9tX0IIOQApBHRcZkxgsoyDpRTywZOBzoshvh0I/x/iP
Pm2Tv7+GRBH/9bCZSjOS90LEPiMO7tyKxy8QGoRTqEACaO95Vrva3PPcq6huMP4Bvx779TBNPopf
V9JKSFTHHQ9quxWtngi1Ob4dGhUC2fbXDJGTq1OS59fA3F10NAJ1eLliuf4g7ty7tPfn1wVoshlO
PVbrU+mfTlSCFMTuePJxNWaIPZCPN4lWMvHnfgsy3GvY7rVGMzHhlVy2JY8g5Y9L0+P5qhvo17bh
Cj+J064aMPUcZ8PV7tw5EAB7YO1VxCUemhOEyvhvFRIeWR7enuYQHSBHp0fTwV4OCUTNhC8bKaqQ
k1LdTbcQA4hjgVVeWC8kiwi5x7Yjb4ySR/bFASRADkUIrUPzTWMBMgOx/Xyyj9cAfjBs0VQl6FN2
ZfVLk/q4Q5XBCJSxZH+aAmtvH4CVM2YdCUpglUkwjR6Q4S8R9S94Odp+7CJ98QqZ5KGiAhdiwM3u
huv3BHhQJn2yfNcIyfBUvmd6Pj97XGpgx/KJdaa5eCeKAQ5SKvRat7FAWwqHXn2nHPF7Q1OcjBku
vV1hELAsQfOeqAjhDe19ds/BbfwPM432Palx5OymXyXx0Qvcn9g82paWjj/B1JfRm7EceIaEQGNY
2EWCouS73NiI2BDFIK0xLpg5Gf4uQV7xbS23rjy8nAkvISK1aaiD31IZ7UZPIw5kQSKpa/LO/XHK
VdCMRs8ZGzq/ICXtwl2ABvZXJFcUT2V6UJlo2avgT2q9sro/3RPY66MIvnX3focWz6xdotXik+x7
SAM8O8A7TG6YkZBHVcBKeAFQGIh5v5Li/rrDvqa2DoYLEECcDs2VteTlKm/MNj8E6ufGx3S5X4O3
NpOe6FvRQWl0VuiZWgax2v8rExtF+fub7toGbZX0WPrsWhTp5ilccPWrwRCf95h3eW4q2gHowZgF
0I5gyM0agg7HG1/o4/PUPXkj1G/LRiQCv3w4oyUprJT+E/M6oAHOIgN0cfasLU+Y4+g/HIa8nyXQ
TMYdj76jm6twbb02DO9SFbNXa5gWmRHLOcA8N9umDP62I11rzEm7HLBlp05boF7vykIo5xP4EGxk
OnA6+jA8+fREhNmzV9PI7HBAAI3ID8uhFN0aoiN7xYZuJ2pfBTFAQTRXe1zCiqG+1fPYf3VhEouC
fGBdNTiHcUBt+kYIgvHs5zxF7mzmlWTPzFhda0EK7zQVePPHH8Ta6NyNyUQzoUdQoyBjtkVHL3FM
FOFYH3SDuWhF4dOya7w4RS4qmIjpTD9zJEDAlSywELX1vEA+GqGK7e/Xp9ewjbrdA2I2yKembDMd
Z+A2WXXb71es8rQpwqxMiWIKZr4SSyrrx0iXYoUNgtdhZuQ/mdYRJdrTwjCn5Sbqpy3UG6VJ2Yhz
TvcZ00yE8lCuB7APbLbcfEV4xsbHz2o5xk5eMYhAfWWFpz1UXmt0agt0bYJu+E9mDa9URtRbnQXc
EpHuJhgjFYD97Pxm71A46pIbMTsgpRr7dsU66yymCkqvhyB7191UMj35VXfDsuhtaqVTJZ+G6koF
nR80P33lrqa/ZPdV7VlehXy3O4PU9ptTujYqJwcc8tW4RG4Z1OnGpeNgVAwDWykhjaZXi9FSP+y2
+37HZUil9+oRschZzbjbMv03KoJxpe9rKCqmeAEL2hqG4VaDpuGA01xrXTOSwvp52MiZWeQLTAMp
uE2LEFU3kWZ9+wMeQ7Eexd8lue11SiOhKZenujPitxh3kD+B+Z9zZf0fD6+svh/p+pPyIRjHY1t8
2EXDkcJ8xF49/n+FGy3pbTmHk58z9SwTygD63GsstPgxoC1yNomlCRbT5Yn04bTGWcRwwA2UelX9
3AoVCG1YaokE6Panah5V1OYwVFTlbQbOLPCMlvtMwpkBBOs4SHD4IylEqI/by8LDiE/WXmNXySCj
opy7mxnXMF88lERQP2JgZx/NIH8wug+Vld9qYmVv0Xdx9Zg44t9NA8Ys/PJh2U23qUStC3y1kxkA
iycgsmw4hnkrzUNjFM84yag18QLTPTMCS+Zc6vDJYmSCKSZT6VmHt3r3jzAWWDmSXCdcfFkm46aa
6SeQJ17V0bYbUSD3L/aQtjSjFpbbvKMWGcAhqTN+Q9Om4Csz1m6dzb+EOSJ7OxE5MVxJh26DVRB2
o+117vH2P4dnFHSp5voN39tGUNNLKz9Ou0Wr+Ub2D88UgAhS0KuvlaenJLv87RmrngZfv5Iw2+xl
Zocq6tgnWRsSzdMMezQA7ywPL0L+lv0MfO4JhdkUP45aEqjzizgdhll59ZCXWZt6OImYuhzt9YA0
ZwzOcYwZdeyBSHUk/IfQm+tWRjhEKcoFvj7DH3Ma31n43P/EWpF5sSbUX0sUO1WE7rXCwzSemcW7
ikGyG8LCuhUxfidZPeEcDpCh1E9nRkXkRoGYsmiGfkChoiPEYsNG8YHkaH492tj6MfFix9QUoKLS
8U93nufC7PtUeaEfUEKRL95IfMM44iqtqY9fGrk3BKZTyoLOy41u/3V4Ld3fJmcmZC/9oBFqwYYj
+nBLFdb03D9p87RH88Rb5VKpnUyWX5D7ltmNbaXEPvb0pWuo1pWNOKSRKDsmaephYmq1Yri2qMTe
MGhTly5yvED2/yFN20nDoaCpcUep+ztIZ0Q0gs1wYY1NpxYhPT3Sw6EI7EMHdIMlt9PK9BqbG47U
aUYjs+ozxfep5KRFMRW6n8saiwlEilRZqwt80UY6mrw4+F3clje4PDoV1WcF+Bu5O+ncwGIv2KBx
VM87dZgZS/7h83ZsHc9/miycQzSvucvVJsMXDpv7nZMdididkgl6dUiz4c7JngrSY7lFvfZfNVBc
zbJz2t1DrFhtz5PuUzgkdjPis+X8be2OF6XqIDpFYNdYPjramPvJ9z3wYAgA8rG6CNoEDq+Y4FMC
/INfxfT9/utz9Gjbh9CtD9BUZv9y3dXYqMyV/cx0b0/5tBX11Fgx6wEiAyJkOk6WFOYXxSJoXNmu
XyTlpmdY8KUSSeNTW0UAIkVH0LA4DN7AnQG7H8Q91U1X1dZ/yGFL19fLSVy8ftjrcbWpl/HzTZnf
bp6Z72NazcfkqbV4QD2cgGE4cApyjhlfS2pEp617MpeAqTwJ5BBfKUvYjM+98QVyDeJ7hI1YycNr
QcFefrJvzsirTbK45YnSCQRtpEQVyST2PADfIgt9vfg7ICKwrB3zKbMIc2RsaRi1am1mMLvfWt96
upFreWduNmyaf61IQL40RGuCvQeHjeZ+nT46Sd4EW3YBPs9sxRN96o19+yC5ZYUPoxTrXEORgvmy
1XQ9+kaEQhBkewlwOVlBoeF+aUVoT1/slkXVmJWLDtiOFxRM7Z28/Faxj+gmiVxr/WmUBsXvPQr/
BNohXSUCrjF0/cmWkcuES58LEZRhehmw10XQWrGxXtNsEsQYfEjyjcOJPGWaiWWbXpNST2ECq2Gn
Y9ENmjZWLBQY52prnpZ1WFRc5R/vA9MmWihF4ZanCOH/OCgJks6eklHwoIjkeottq66A9+5rajht
vbBtyLuoPX+hIYPy0xIKQwfp+MnPCui9FcwZkN3Zyl8na7RPWTc25SzqLFr6L/tcuTdfXm1439cg
QCpsdS9/vhol2XnFSf5hIvMelCtpI++x0GMl06ZigDgka0rJECoAskjCK6FcMX+pWQxfGXkGvYIu
UIXQsQoQGq1PTD0jkZkL3ZtSpV19zy2PJ74TNnZ9dI18Y2vOLUoKALDQm5PqPmkPBznsJTTJntZP
YwL0XhUNWhSTriDbFF4nEDxPO0it/cUo9h3/5I2QbfLI0J1MwTSwZg0SWMt+MunqEsBy1a7Y8iI3
+S4/yCDs6fGn5WmJjGPpQNiHVveOQSe5THjLDrymQsbP4YsXIxGjCOpoRDlXsYanBGmFfy0+yFjk
OHTFBbZlIoHkKPjCZgTcylqJiSyhUx56RwqqvY12e1haZKCCy2SlRuTN9O2vL7+EHv/x7WAIbayV
6xyC+mmQCODczaV107gVejPUAuT1YiNZBbl+sr9PC9U6ea1YxmiPwmA7AbxLBFm3rp0QffJwlUer
8Ix+GqJWNsVkMLcxEJduILfZ7ycrPCsIIc83vEfkHlFoTClOOck7A7YX0T1LmV+WKsEhkIXuqJpx
xhkHvHIifMB+ITcIo3MR4j0KvZpGT1fq/rsdebUXoyxsTRzHSfa/hNkGmCxbiFWb2iNpa7A6MRwi
xth9I0lii+GeEDFCsWdswcixJgVACyMCqvjQKTHLiABWx9nwaPLLMRIzrAPcxGYWXLogFWQrQpou
Lm8GCqtILkqrw+JALdqv5NTsFTFkDsZjC5qa6fbt7Bz8SBUx7aIXg16S2uJ3EamPrTmZ2hAhVxC7
01FbvzwyiQkZGOZfUeI8kD/9gKdkZaoZbAH+inBGWnCfau6X3SeZ9t/obkcZ3grI0HUUIca1+4YW
Xc8VFIv45cT0pPSTF1CPfDmTpSE6gtMe2+S21nOUQVdqfzfGVIQ3S0Oq0gTr1pA8Wy4kBlYB9qLQ
5JzVM8GeDCQiI44N4cT1Bkdy/6OlRxrM0bRBkYf+Pz24RV5Ijjd4WcenYwSabXbKqdSNM2W4/oY+
AgK3BFPmzL9feB0HK/7yKI72C73rf+wgt5McbcDPYjXcRDDDLXKwsMWSoB2om3Kd+kOrZJ/FKWG7
FrCsES0MQ4u9AXJTd4+rzRrHas90a7N57B2yEyJJsEh1l52USop9DruKQvxl6qwr4LiGeXn9cHVT
xcffd6YjlPfY07ar/Sq4gtIKWPXt/te4i7205pk6bSiLf4H6Qrvm4QVnxuagk9MXa4XzisgZNdQZ
sN80WIX8Km8uwOo44AgSfEGKIzWw2S4PqlEBCOdINiu1dNfQw5KsRZsRbE1EgO5GY6ldmRiD0VO9
72A23TsS0I7Gj2f1ZjfY3VP+dPpgBer70lTZb1IK+xbWh++aq1UlzEkQo+tG2FwuWMNxnjtwrelW
n8odoFkPfiQkBNrsCssGBLJXyIe2kxEcvXCC/k9rvJAqM72osEUDW+7Ocll9km/nmeFRgPNC3Pma
zuzUSvJPIsTlQ0NLykmTL8KTE8M5C+MCRSNU99qvgVXlF9Ta9dqFCzyZvbYfyJ2kRhpzqERRz/yJ
8P8WTJPBLj2Sr1NbLRWYn59ANMD7BM/01SqhXHRPEhmu1LXCh4XQvv1LXvCfrZ3Nc3/u6a04vsWk
J2tGck7j1gxSbTgxaAGdEupkXOu1r6fWcn/f0K8UiTGG/SGTezJMAms7VykADTgf2TYyffbfjcif
fDS7VrtI8oRPj9B1rZxvc+h3xgpUXEybaEkXHyxlFR3mC7LYlHUV19qoLK8azb9AAMlzPMKrrqDz
wrNFP0XjZgj7BmdbJH9iDZEkQ2pmWUoYgBcFlsLQCAZPWjjIRs1+Vn1cIm7k9VnKf0QqD45POg8e
KceMk0qmLbvu/3DSoC9IBZS38b7UcRZWvqFNh4VsiRaPDsorf1YuhAVMhMbhiYBx2I2WFL/tnXeG
AieDZgyHTYPKFg6i2wwmJwqYOwWXnLtoB2Bon0zJuehCWNjjbt8m2jCHmmVPEV8A
`protect end_protected
