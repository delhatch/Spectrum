-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OMhad1BZhDNpjCs2Vlz799lrF2gLwRCb6galnmKNVYaR19RufzXSs4PREUlwW2UoCo2WZM8RTlyh
Y1TcaMGy50LxpS5hMaMUvgI40/nNrRkpx6tq3zMs+jxF0t7Id/abD1YNTYrf7p5sgTq+Ppn3Y05z
4jV6UyozYXGjNYRp0RLqpRSlp6w8Tn6YlBbPFHaFQ6QGH9gHyaZfOH9WSg7SuHMLgOHNzS/KasjX
700UKnu9ewFTBG8SKtWOux7tcdUyh/VEFy0Lc+jJaRn6hiWDBm409xMUsIenG8ovOs/y4+ic4bI5
PKSWuiMyID9hVgucU1aMKZUTuWEpOFD9jXwqYg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
DepfBWAK+nNh6bVLZYGeI/FjouwSCHG4wfegaUr/d6VhPqFEuHsXy2aYcSJZzo4YEFr7kxuWlQOM
voq4vIDqRzHuLteqC/t3fa8SxuSo5w/q8KVlWwCfimAEFsIKJ6S+LH7UGaIRsy5n9O+yHMhBU7yP
tIRJgMK5g38n3tQzSjFtuCvB6PIokK8Ildhye1JmhyZmO5Etsoxa9wiblM7ebmoDWb6i2O0UFJQ2
dlhp/r5BMVvZN1vpe4tdoiqGgBfjvUMtpbyXBkyxpkh6ykbNMJDRUZkOfyfRi5/+qU0spfPHjPIP
LHctW1zWf3QxInlKZbt6xWQHxPF7SM2W5DSwbtUwcaCUd2t67NJFqqHRGJpSuOqBpi2rvZzgoVWl
BfMMw+x8yeMD+giqxEXLWgFB69mkr6a4iIKva4tYyUViDst6FhHSaFOprkWWXuQAaET1+lmR7rXr
PJje38qqLhuxAwGRej4aILkwhcipgVLJCEBcyxo4oaMzPvFGX8Wyjyyn80FSCtgOPeXWvRvwQBo8
eSfgd/NnyWJolIWzGQcDwWV3zjkVSdMuUochOkfwZ/ilwJdkVu+JvReXLmgKfF6wEaBUxQmOmIRi
tUVDnwiEHMGHbNroEhwaddOx29Rh9As/OGylDeJjAQ00MjnQoea/VuGFDvaI1iw34BSQv26ZbSpc
XD/VBiyrvK6jZR+UWwG0f7JB3LPY1UDOADOivc+t6GF4uk6ctBqSrerUWpACT4MxuR2CdRFhmfvG
K8z6ZA4puinbDvD+2N4OOaVfZ7jth4XiVbbyPgLWcJjlqZvmHKqMl/32Gc9ysy64wQDA9jTlzMAz
H/oV0gyjGGEXLgB3Hjg/+DgoB5gCdGaqWZ3N90hbpvnpBjyqkcQ04elM6ImgPlTBQWO+kdwVnbwE
lsJHP01cPLEj1AcP2q2BgBisp54Wrc72kRfe+yLw7f4+kz0FoIRbK6383lXKLJ100JFepgYlwM7G
rCIsJD+GBys8z2vD9qhS5QCOi0+odcD2IWvDazm8LYOrnYvzjySzpHz1rKJr4gJzmHdMzk47kgDa
ubhNTkTOjPkbQsSOEENfFgo+trvtU6krcv3onOR6zH5vzv6AKZIWLCflRhCvFr1L3zot26Gu9ErI
aC520ULp0RN239U+kWEcPZKFZTOOikB66E+JsyTZgFRh34TFMxvwOvg6Aq3abXYnKA41WUcidH47
ub3xw7eHJ7ZOpzh2IBMq5bSQKL/a+6BzElAiPIlqrGPQ1UbZ3XKS+7SMXXx6PraCf6hI43vIzXhG
l57V0t64bV9RpAFNoyFnuCTv95p+Bg9B9MGEmj/D+fgNkK0RcHKQvnG4B0D877wAeBec4+6IZ+Y2
ZOtCPlhuMR3Oq1hFzIMVQAm83gB76BZYU2zqdMusnYLOFHKNZSW993K0+Xaa0OEgpUDSdQC95ulk
/vLANG9Y6ewi1wg+eikFHGM5GFsharyMOXhBQFnFuMpAKPa0xWuzrdSFuVmIgtuXShYPxw1qViLW
5pd38gAHXkam88TmbYQpRHbi5jIXKs1dtMJuRtQyHj9HCWFQaAxvq1ckq5wZ02ikDcitLmdGEn4p
iGj/r1L+6y6qQyiPdeDW9Ok/L7cjBEES8DiAcCxS+7l+TVpuQQ+3UVrXIO/c929TYaz8JwzJo/6b
P9GQDZNqzUeMdFYgYnx+4y7Fu3XJmz8xB0u/VVueBoODGaEIpAe0xXdhXPTlQAUY13mJCGRM4rNM
0smx1pnE/uNfpGlQCPLteS/DUqyMSRm/w0JPLRna6LIbk8BYQfhvh7V791nu3/sVXSy7ZKKa8lOn
e0i8WuJCOgOGw3mskQDpYAExDYiRDAeYdigtzQyF9L/JGzW15VUQAtifHfNRS86WwBgU1tTF/9Ec
GhrE904zF501/IBtqzgiusrMULCdTNNF3qBuBW3CTr6AJWuxx+BkZXcBowX/u0WqkquZRbcImvwV
byJYsPWKkL952L3bhM2DFc9DHdH44hUYCZIfLDfl0WDSLMW8EN8dLjFZzQEmI/luMlcs8OjNkC6d
2+oGhGoBuV6n6aAJFnANR0b0ZKelWaBiUd3g5Aq2MJkEQI2eykHuoGbgV6pm/k5oNGpRfemCx6uL
cFnaIeWklcFayatBHq77FODFeSWtvUkAl+MarcBKP2+XusgmYS9YNflk3oyjQ6ihiTzWhgNQUbFu
r9tzMqxn0QnGDwH8pxDOjKREGB1Y2DrFQ9df85Yerv9p0e12P81gPmdUJI7DsdRbKXaSlQtZeegB
2QA8arF/SK5qAG0SR98VGBZdlqiEWb4HDzeeMeoTcFZqW9kDdg0oIHJu/doUWE+BG+M3oA35Tkm+
4eBUvcmGnZPCnHO46FORfNtGnL+JHMws1sFfoUoINa2aKNUcmt2f+L7flxMvbi+9VQhTM/+RxDEV
NwoHM1DUtLHSIzUSyqgc+H7KIQIbhH1yYs2wewaQ69/4jpkIzqXx4i1IPdn26BzOj4Jww3weZOD3
zDBP6gM1Oe3micaV9ymhynDkkFTtxiG0A7dui3f4jdt3K651ftXeGrCBK8vNFWa64wtrDw1q8/KW
WksNIcnF8Pa+shS1FOPgl5h450cLnVuaq73qxMRYTqle7GpGdlWQixV1wsPsut4XDVq7nn/TosUG
jSwf/oe62r0V0lvgMKQl6pyFKNTnR11O7ie4bNhvSM7zjKxIFnUNpa83+/T7KsxYnZbFB/jJUtWf
dprxmaNKzgy2QwfxAcRMfzJi0ITMe8vU7ApegcWwgARVBfz2R5v7/i7yqbn6SzrFZ/8Qgh1Lsq2W
2rOXn18Vv1Pl8ITqd4LVrsl00J6CyCa9TFwehEkIsRsd7nyft+wrsOYpV78Lyh1XSKFIuLDFJ3nc
hdMIhn7VlqN1Bzthv1UsxFpWJZu/HqeiBgVEXtTJwhmMvwfzbytJOKlYswcnE4KjY3EXLImlDR8T
uUEkla5JlgohH0U8F932xemYtgf9hxPU8Kweoyqerzy8nqoQzLiVnX5sM65Fqi03zenkFM4/jCF3
Qhr714iQbP4EIJpS/HMa9P7L/bi3vW5qGIioyyFs+Z3lzdBRmiGuVDWhqmDrqyKKyeeZv1EnZnuv
51rQgW0pYG+OkzXp42SY4SU/lnx/Vz0+khRe+SqI3xRdIhP2ImgkO5ELFz1bOGBzrLLi0clkAenJ
Xyu+jVSEVSBpE/h/Qk5okU5TDF5+5B+EBmc0klW2A7JtJO5sUccGMEJTXIzhl71Gu/cE0WbNJCcG
Y4KTCpkXIz4t/eC3OFLyqPd1ZqpuQehRxq+mT8N0xwIayWnEPyL4Q2bLwYxtYkM1K+aNfIwaTBx7
0/yNrc0jNB+1b/IfxBkv8MJMhdT+FeWoWmDYHfbGF5Z/7FgI8Xpwp5GZG5xkjJeekK8Cso/vNyzc
8mMxFC1NQs9d/5CtXX5zLPLAGYMHdKx144XZXORFSvPPAESTku4N5GAPTpyezaw/7yRM792YpXB9
4wP2OeVeh5aZplgPMAYlSB+DV5Ofv2qGCRO9VGD2fXVA+42+dqOjU/jrfRa2cCGwS+PYkuBxQU9o
JASPXifSvNzhqFLglbPhqV3rZQTRw/0b8TppsHpI/CJ4o0tWn5p/s9ffEL/6biuD/ZT+QiX0mDiO
wrtAdmeHj9W9aGjXqie9YRYdn9/FrOhFfOBh6F04sQdBzxv4qdETJ6rwR4K/WTa96Ib20HnzCH8/
IYa/l9L/QoRiMRb7FmvrCKxvzHYqzl6O9Ls8F9wBzXKcwBrBow/Sh1T6VEp9Sh+ukQnJXgYosqoV
BXomWoRK6XF+34b942B4XolDQvh8SISSBrwlvvI/r+nIM9VO2ApBXAfDRxXJO/6GnBr+vyrXVdlA
x6KC0AsIG/fq+nyI81lKFvyJn5yR+381zfB2AGi2lIT6c8N1uiy2b9JIAwKgHqoUKt1IMv7k0G+a
bsfZaCW/1HxaC6S0pPv6gst/xtkmSUzOIvmRD378CkraFrKhs2d5YEy/NV53C0AcI9cLNGupUoq6
+nlfQTGDh7IJ5t5sKyPMLaTslPJ2vlbOe0f1TTMYgjUC+s5srVxxW7eu1wHx2nLIhcXjhLxME3pO
yiSKa/5MC31lpZuRHNrtBmMD1ilfiHXmu09BD5D45rY8N0QUYfi/V2e6AfEfhFTARI3Rvty/dJu4
eUmMXwDZU8hJDPc1vJaIRzYAE5r611AL8OU+TQwPp4BVMaVzzV9yu3dYrc1p8eZ0Fk2PNfXUsZW8
ljSfS6jGkNbe/4VOhLNVsGLnxzhm5FWvRtrJfsNqknj3aTP3yk1TeKKVdmx4ELEPolen2vJHIk0u
FVW72aWp53jYOFBQK8+ZnNRlnrMaDib2vVhcUNa1rTHU9j0L0q0vc98wzzOAxpZ1CnPVAHkFAiXf
AMdGcPl/G7p1e5L0/3o24Mz1a7MxiNdOiCeySLsjQVZbP++NEOg0NPHwuhD32W+2Cu62ndVH4hoI
YJLbiomgDsvogbIfb0NzoITW1jsl+zeVTuAr5W6BixRzZd1O5ntVpGWG+slmJ0kfvV8S1QaTnFsT
DFoyoS/v9xLmvn7jYDhLOFA9Vx67s4XzakdcXd2YZZm1WN9MXi8VWOBRdFwN8PphpMogTEO9BGrO
bglfavQNDfuE1J3ujXZrxmJlFhzCuBhF/4D4a3jGbVkJHdOEqmjOxacOFV8DHy5/gYrrSd9iGyLx
TOxHMDRWzfkqeMJyUl1YV63JQAx2xq3Qfln4tmSe/Ivy2s7gEaAm4H6ebUTMOg8GPUEgNVaR0jXD
/GQl9GsL0LtzGLvY6fFUmAywHClL5/aUdS0BsLJLVSFPRpbNGQlXz07OIaZtbwqh0avF71b3Snoe
r6WkxmeWuYrQfOW5pFvFSAyR2R5uHzcREQmU40rmXPwlvSrM/zwXw0J4ge3QPrmJdChjcQCa5PNr
KOVhgLUwOZAUwno9iSy3mDDwHhJQ7uZ0PatJoDo1kcIewX0AqyJWwLmgl1rlqDbQxrXqWE2UNiqa
85pJD8xhdum58yN7c+FkWMcGecbzrbDmILmiIVhEUflpQRyfjUx1EN6kdnv1lDf/GTAZwC5IBR0g
z05l/yoPzVlAPjnnA7RKpXIk32hghfv+cNf5SkIuQB+B5z1FrY2rCWNQ9smV4qzwCwl26nhOKWKc
iIdbjxGBcs2R7veTIek5ohVNccjjwCSnqCGzpSxgaZqW58AeaCqDz/Md1qzkafewCREiEbpVx+yX
HjlnGSM1B7cFgrpeSa/K8YT+CUbjANAYHU3eONAS/of3S18M0qB4rpBlq7eXhRLZ2ozr9UNYd13h
xqd3Tkqg/xxDf6Lc3z2hgR+iHqENCO+Jw5xaY1Y7pHyxnY72JswSEJKg/C1FOU8sPnZQEzuO+3H8
uXPbYixFuMAh946vpXGV2kG5rUUmfe565/kAQCCvkqjc4NMi7M/HlqpWRWNuglbOEg6/DrNijbqg
P9+1peyikXxGLzQ3Ykm3sZJ/lZhz6CGzopmMGiRGVmAiW8lpjD6QNHa9anAstYKGuZo7+defd5Qk
zgol+NG5cnC5/LdgGOFnTMywHlmDjR5gOowD7+63Bv5ZLDY+OqKyd0cUC7QnMAyZK2SrXnCeI6Px
QrjPzLwTGS4XvzREiuB6gVpMauEtfBxC3vaW+nMn5TkE6K4DmN1uAL2ua0vHdX6P/89YCFsOmZSB
bXrLY8Pca9eqEjR/mFsWuw7XdFVPpYSqB7SNQbaHmN3y9SN3rm8kn9kS5uNGcFsDnvbf+0Jp7sjT
0sc0XMZe/R+8FQywlh3wQ30DmrDHE+phIevZpAU3mWpiqHtm/Tjyir5RaMHLOK6uJtVvsQeywPXd
UrNyg59/8TjhqKooxSvRF6loCumHeDsrA/9Wa4Y1PD4c7TDYpDzUFHCiZXlL2dQbzeXC9UKNKKcl
eScnjN3QKHNNCOd2qlHEf3PsjwxJxKVqiIZbIDaPWLfC6Ob0rPHvdCXLMbmnuBy4wMKSu2xqsCcK
6G306GpNc6Bi6pRWMswUtlGn4sljVAKwAdLFtjU+9u21Bq7zhPbOYnq/LR3SIgiZMBTL+XysRtKr
NQ58gU6esfdGZgwEv8bgzy/aExZogLVFGZtBvyD2S+NnHKbx3h2IQQC/BY1dIAhD6pxK7nEWUKqB
7MJYRKVWqam6fAyLEkunmvN5NbFGV/5tGEsZnbCM5yhgzYopQKx1AOOLnRMdjpHMw4CGmCtvuNje
4PBDp587PZiloMpM8lU6eq1T6BOgzpxokgg6AeQ3Ct3vFqafthmqBoEmU7ykl7aAoYXt8uYHpBRO
TfB3e8EviZcZ+ZRF5Cfm6FiRvLJIX1LnlmEFlMzMPQvrQLVkJgfyGvPpXNlGAGXgKjJ1Mm9WqNJ2
4WnTtFIicmOXUMcxs9dKNOo/GmCwLnOG+qWOt9tscXCt/GoxyFO9jYi0f4KmG2+M6mM04XERK5/V
uDWmUO1zkZFOta1rN7aI09IJY5Szl+g+QOmd1GP17uG/DmYs3qcvrK505GMhMotMHtpBuQZIHChf
dvi4KsSI8cygxABU0l/MZ7lrzHDgHbqG6heR5fUlMgup6iPRlEOQy10IXy0SoPV73zgpWr5qbmS/
HQxQVZErHrMWu6PhNQZsBmijUwEhgOT5fn9rlEltdovte6vGHHkzIpDPzzpFsSfOrcQpB9nz5rj0
UQnkcICfdNh0+DEh9a07Fui/sV3efpJMjMG0N3LUG0/cPkHwEGK5CbTy+7l6SObIPaVY/vvkOUeE
o8SHOSX8aADXPsCE4NrOZPjuXCTxZFoI00qGSz7Jlqx1XMcTqrEAcPeLQb3RayfoH70BGxRsBfzZ
qGaeHJFecRlXG9ietZ32s45024bDF7VLimeXzuRHZrec+++AyQrqUquaTxZComEAzG0GDw6DR/6E
0YvJPyo24vZnEFrVGG/J1amnEaMiG9hljvnt4FYTgBEdnJrdv2JDfVSrcX8fzLR+wBZybzFYVX36
DHKZDWG1JiyUTGHkEj71TlYqiJHhonH50L3hr39q7TumKI37OT8DDIFFtJzrwM9PSr0oJ+usqDvv
Z9wO1u8+lrZhG00I/is1NNIUYl0IxJZRvgjejwbfgHTW2LmwMQzh457J9YYdZYSp8BktBAF1sR0B
eUZh9nXUWbXtbzoBxHQ49BR/Il9ii2Q9sURmHXzihzafQTP2LAx2y9ufUPWHya2Y2BCSEAvAncyM
dJhyCJSQ4YUZ4co74ZmfD/j7OAwBc+yr+b9NFEkuigD0M4epeVL8r85+zNKiHemoeNyG4zXJYz9r
E3afgD4r4qxEDscwkfU08bBbsZ6LQqDu0kjth4fylmMEYImPr3qBrFMe3qGyOLp+9jPRPGM3oMh3
gVOUSP4Hx2dzHYB9qClRgeDgMyeUxxkkI9EqYOqIwT1dn6Ta8+Ri2Wj56njBOX5EaUkiguEXZrnl
0PLgbsQ8YRSxppghTi5tnG0S8k7XnP+dTZql8L83miSXKgdzBt1AP8wGQIJ5fJEzKZUvg/NNT0lI
nhW4DeAdEWt1CxagFmRxnFSYYoqutVq1xl+ZEJvi+/gVHmnPQraTGeIO8u68CizvIjPd8Y78Myyw
2fd+892LSnVXq0Av/lqfOy1J2qLbnjGk+bfEwLxHTYthzYFm3/6qlLhN+wz1RmiqxxUh4xp4f5Tb
/eMQf1mvPBYWK9Lz9f2w0pIhhovSgkbjI0gX+taG+0O4fmRMkn2BeGENa6gmyk0R8DjiH+mFhTa+
hJhHAvKNHOjCAK9czwH/gF5D3TzWMNNtDl+RZ+giSeZ0RxXHKLkRgNxtf1SuDKpOr00KHKOiX3GX
zI+jgwDVxn1YQx1ELoPZBwClkDjCnE5fy+Y7eotphNvWagoK3miWyeRZTvhtzdL/+iSL8qNgnPUt
POzg+l+aO/WK8A0YfYw9zEWPNJhNPnkyJPqhtAtGM5Te5shYkKYIeDNbEE7bmTB319F/gzWiwB1i
sGxS7xD2WQmgA9nKMGvQAs4MEHs65Kv88LBSKw98/fjNycZnEGOfdI6LU5ppshl4286IyAyF4cBp
n1054mYfjTCJUOtKnCUgKmBjPJnVTXVJT3I9cYSwHOV3XYVVO57RaUSIstMcjvIBLTo00cnR6TGe
KcMsBx0YNC0zz3lXGppt5nDGNOF6xoa5gntT9sByw64LmgFD0CP4Tsue0Q+z0vG7+TcXzD4jaBTX
zbp6rMQU03MN4KCf7lIvfdPg9DrJdAJybYGRbXQdLT/uYHU7aop3KNeZvJ3X81uTlbWtHaoB7L5X
KYD5CQoI1T9hgoGypZtg0bybujWDw65xxx/SXX0OCsOpzsNaUpQDzCbQMljUVepzBItifpMtebgj
n3CGl9sbVD86H0vrZmIUUVYMLkHGY4xPsDh4V8tF6XemQv2cjN5Ryzyikc1KAUDl6XCqHOLgKDul
+r7uus/BuYTiF0E8171+917rtpSWYT7UH+wFWfrpOFsS78t0dEhq/ZCI0ncptCCH1EWULnnv3PQG
McBYPgRhSYhxTd7NNLdmG8ZPzURxHUcYPOshI9j3BvM+YI7oj5HKYZXP6UHmqrn668ynS2td/p8V
++Lc3Waea2FJLxWUMUNBWWFN7qyDirtL4M2LWPkyV82aB6Y0YOfFizTNwZgNecIu9pT4Stltk1EX
QJZ867SebODTye/P6eR6IijF4jqdJSqW0Ze/WM1AZfLpG83pWzwl2FEOlmwjTUXhVR0XI8i0HC17
cP0W5q/LD2z2ka4NKxBfwZ0yJVGmBdqagOW6pTV8bHr6hcW6+jAPiA0U3gWuYMx9Kbdx+nLp3tIT
vAML2GOYUkeVTnYse6l5i3HLhDhMNA3sA5wG7L8SEHhmv7K0nAleApm0L8RdIWgB0h+DZt+6/s6w
F3PAD6V1F6nAOkO4oIIfNgKnu72RT4X5EvvChw8Iy6Vt7M/a+IcTUr98Z1sKrtSA8ABaLusf45VT
fTcJ6jxB4gAhLPM/cEHM8abaocD5hg613+kBRILb9JLp3qQG1aIkRUvwE74n1MDW+8jDqMz4ZY5D
lLfsyefRSWA+uwHDfU8mgLDWI39E+pOpgZZzY2u1u7MniwQZ9UzajOj6EviuaVj5iRz6Aqv4cYpA
h7o6Xt1iC2/sHEN9ObbzcXQn0sLOuRe82K8+cG+xreeNEJKRxSm4FpRs88qBrM1rL+8jNvNOYCQe
0aZ4bTzNb9PouL5/ptGxcG3JOp2QkvB3ZMMGrSEy2dI7JNZ6vzVQ827o4fUgfnMJMKPOAFR3VphB
7lKwxOSlKKZAyPXGNXDIReLjaEWKIc8rP+OySBPocXyHhTdTdRbwsNWD2CKHpGq/CtrDHJDyglzP
zQRWDykXH9gQGNiof0u3G7EZFn++a7pEt37Y9sALlO9Qgo8sy/PJhdu5miAsGHS0ewyR4BuBn62C
C+6ZleQ4mVj6u/62CPq+HgDQRJXRLLCxcMkho+kxbClIHKuQF3LeA6o+WXTw0jw1m30g7T51qHoa
uJuVGAhUSjPqPTeQLZYZaZCGy0uLjzJQ6YYYAuLEqA5+0PE6PoKv9eVFXVrQ0PymNO/NNma97Ai1
zZBGDdNgGfWTwbRZAF6g/I1faTBfRtDfDKIdOtQrEyZNvsZ6F8C6zHiOf1EPQqRNcQ6kX6P//zus
HzBnidEs/XXiAtbSkTWpFVImMaGn1HkXvJhRGI+yEaC/ALi9DGwHTMmEMbeopWqdjqpDb7XgzR1h
qK+rYRRmYbdxcnxqJOXikKVVob4i598TdhC6I5K48uH0lnbQZubrE/XQ11EEfxMQEk5pwON0obXj
rLoqkKCgcYAGBD61Hmy81O5V6fO+njTtz0voJtNdJIDmYPLG9cGPqXxAFZE/I5q016EJ2hOzbKXT
IplCaf0eZlCaQWuL+rVhS2GxrFgVaV4nttgGwnUNSn/CA2EwagVbP7zS9awBQHYDA31grVP2y2yj
NoyQZIfteTVok+WuhPRQKZ+lUKjFKpwcSsx5IG7bucSvDH9pY8x3xxYMQ1/Pqx8szjI3uW+tT0yz
VedZX971g5lM7BaQ/ILG3lBtn/JRGuIfnom99DwR+Ja/8uVsiW06CTQLMx36abca2Oa94LY3m4fT
908KbxBGxGa4vqbXNyyzeRJVZKfG9eZfJtCKqBmJIjL6XBLhlnT+DnXfUiU6XAIjP4aG5rMyvHdX
eTpaI3ObJq5LQyw6R87kJd7b44gOKf5Gkat8ze6nk35benezBg7aH7stNVjKIRSlf1VU2B0wYBWh
ulSfP9jxDAoO2c/CtFPwBxfR6lDHZLxPYWtynluBt7/gaIOjIU7aOtB/k/HQ2arFMsG2yHan1W2E
R3MKX5VStzSJobm/8Kt1a5PuWK+hTvVV62XERCtRhDuO3UAGeqdsn+64N5YqY6NAa6S7rIGk2Mtq
Su1/Wpv2q2DJ7lOdFkA/DA/Nj16xWmjcY9dx4d07jutyS7d9RYBC9jAmi8RlS+8Wb01mlcWZnD7U
DDTyBcK5qJywnUNa7v+xbry8UToei5hwVZt8u1YJCddqR2dIGeI/cG9QFoXQpi2tjdO/9NnHOfN+
CkhI3C92r5V9MdELIzSYMj+h7+mI/EgrMDrhXOHJsJabMtmPwJR603aCvSARzfEjFez8C+ryNA8t
SUjDxhzjRy8L+R1enBapXoL5poNs4qkQBWSysG6sVE+pC1dCYNJw0+y2/wsM7dLHl3VeftZ8vnP+
lb5O8dh1v3XkrZrfqQ6cYnAH/nr5z7U2LoXF/pNT5bSr6I7+2hiimjVoal/bLj2qS2LW9FeMQtwK
orS363G/xoa0xo4QTvRQ9qNzh3KjNF8m3oRpDl4RsUljA+N5aFl1fUVyvKDXKe9SuAJAtIsHDC4o
ElYVgr6/N0u9EEpRO/vDMc2JFc5FnuQoGn+scHPYc5qbGdMqfPDpaSh8JrD3D0j2VnOlvo34Zqov
ivnG3SYDMIgGGFTd42IXuV+mGdT4tFnRQwJh3rh35Z+GMAlijMgeoP8S8+pt80z3C1/o7t3MiiyI
MaCsIvw/idObePz+wy/5XvlM0ndJ+F1g3bEC9X90G/d0WHCxUc684Ssk7CQyJzuYUSuFBOZw+6HC
4DYxvY2wCttomWXIoDbSl+Sz+3XZrZ/2AZt69seZTMJkn80P2vY3xvnHAgIjvXaBx2cv7EQgOzY3
FdHlTWeI5uT7hU19DdiDVxmGw2huitE4zEnz/4Ry/wERTGGfSefu4OHBsJYG9qnjAeJfcePmeGAl
KU/QjHRTtGcTNZvA2OITEa0H7WYVF3P7lgy1JroYBnGoq3xm1Q6ErBvs1iHB+AYWomQj1ToTn79x
hkSboMOXYH6bii4GrKd1dMoHl05+JCK60ChvIPz9f1OnBPc5c5zZDPwqFwurwG5spfiw100Q9jdQ
oY+exEhWbeTsdMI91rHRDEhyj/CIby1l4Y1tZQPEbIFG10B7oizJszqPs3G9Kvffa6p8iFUvMjc2
VAYJq2iYIBOrjD5OMyDZzvKtHQ83ZQFbWrGsB5efxHwVsQe7ZnzqMp5icOxFqgemm+ZIMqg1YF06
OkmV3yOt2Qtd6bntfGTx8wRUizojmlV9lFlo4hv8U2Zt+ZNovDOF5MuLbhmkYuAPGr1Icr+VN6J1
dKm0o51WScZEUQxplaTWcTOJOtsE8vnWdEXIJPpXDOznGWE1foo2620a6kqpMr0JIcfInLsrWBAg
nEAJBuWakQRJ5vAlkt3z7t1EdZSFWKnRSNgX/1jTFbaLSNyKRvSnJQuvCV10ZDWqtWyxCvAl68d9
/GAxeKIwBeYUN+PEWU+238YLM6IyEMmX0IKHgeVK62ousHCUloTtVSHCwJd9rAxGZ/cVDmoCsLcr
YaaKvkxN+pmGjvNtKkCzOv15uvvKqCGO5gBiWIHTi8skFEI94Lio2TtRaLb5eNEF4qgEZBXJAUPP
gMl/fAHG8wWygydyHqJ3QCTJ7m1VdQfTfXf3pCE4ItHbpqU9w4JxXhZcPsCUdwwVjhyUQ/NNjSUX
sup01n5MBt2JrQm0zMdXm2+wa35DkaLS/aE6du8MI2Df4y9rLy848P/0GlxED5XNwdkch5vtguVE
1STh3dXiNTFR1p+2THK95s5C7sdcAeEfwTxkm3axuxBK5zLbbqVVYx0e6Vn4vxe6h52NX3EwJ5yg
vCwYY791b+gtOLyBxwqKaYkFF284wrs0XmPvDrGWs//BXsM7wUvQuWXH/r8NSBn3lf4wvzK59YiU
IvqcT9CmQR1ZIG6OJAYPmS0f4boefAb5PGSQSEi5mDQff6UchSsEr4dzMXp0wlIxAMHOS3KobE95
NNIjJyZGYEvUTXmPZ6XWzbkLO9EPB1fkYDlochGKmrJu0lWtx6ExYvMRI0F82sL66QMc4NFv6Qmo
2YdaNF+BmjNNq2XyLMDWkNbkzqUMNz2zKyBGLbKAuXil1NLkBGqpV+bJrHO665foZEcM26lj3zw3
twPtSQgMgv6mx2Dm/gdbhsZqbmb6wKWwMlPIG4zeJyYvtxzZlEQKjfY/u5pnscHZ8+urdGCvutM4
9wLnxB6/Cc/Vt1RSeQxbk4Ti6yckJ10N2Kg2nv4sX9pOYwv+MXemytKt5wX4lwKzFpwbvCJY+vrd
TsaLn12ur9PHIVNXQhDpBLC7bjydLnGhXKzJKIV/EidWRNEdV1xLv+hzmkjaJPiiEBj4sfiY7xfk
Bq1Z9vyEg0xGKZDU9NMcci8gldilqeZJ4PkcWr3KmzrRS+3xbsGI2MKktr8SyC9tX/Nw53aVTqDp
Dr9/mEQvXMb4P/P9t1tT+O7q/7VoIg2OnP0xNfB5Gs0UO7yrMiFmE3zOE2kRnmsM5jKxLmIIJPNJ
yNdFehHxB1FONAiUUhM9kDqtLBSbj9r1yDem5ITlx8msVmOcBs1iak1Lx7AtqAEnT3LZyEsZRbzO
bb+GoGGpQQIuQxWhZsFkVtTncSEyWlWOlBIHsMFTkqbmq4E2269LXgGvBoijRf5eNFhDbTOME1ju
FrqXAt1V4Jg/7j4yBZr+YF75IMMxiXvErdD/BrBZHebNOnLohcOgUrgTpx5bIk5+ZdhMYsH4kKSU
XByZKQhSNaBlg+bCvNuDWrRJ+q9onog4C2enAgj+2RHvUBAlHCuwWSgib4rdLVRjwvV8tTvhsZ3k
CNZxz4SihzvonMqPcwRsFNExYn1eoDX/E2D0siUYH4X/rfF59P7m7zzsxg/GeksW/9hvHRJsOl/u
z7gBZezdMsFIOrztG9zAjP0uQrPiSXt/Jh6490kIOHdmMeQaAWbwJKooPtB17Tf/5/KWpiqXO+Pe
dlUdptlFOEdPDftmPv2JTL//E4dljZz/EeFXbGfbnZFnRAvpYF9e+yADdHaCVfkIHodtm8xkw+mu
eqpdzKhAcDMYbgv40PShdMJulezB/rxuZ1pdWi8/S7mtnGuV7FVc5Ux7TKCHoSfFiYI1jNjXmaCD
xJMZrxyZUX9N2L4UddO01iYzG4HRJ7GgAW3cBU0MT/OhESkF8n9zdEpXtKeo0Q/BYDENtqEbq5ZQ
KTvRwX6HY1C0sUNcPOuuTyKEytVfjg0LSnosfr7Q2TY8cxGCk3+9nlddwlvklurhN3vtdHtTG5du
qv/Jk/m0d7wlU4MCZIU7odLLi+2dnPZ5Ko2H5BVoQyysEZdont7elj8DrGuF8jtv1jHr3KWI9yNt
IeU3DQM3ct2cX74Lj49hwr2fZRo3TpYjvZNJq/yIFiQed+hWZSAJInJn5qU53NABCi9zLh8SQz6B
OGxtcx47osYcWvMpnwHhxb42pZRRKJ6Bm8DvKAVH9NT3juEo9tWVmazjgC1YuyICtTP2+YQfjyFf
v+qWhPfMPBL/EN//uxBEV6YVBCpxT4hf5XtuyvtcM0ZZjC174L2dHvIa5IpWB+e6r6+T91oxqFeG
rmvYG8Qp2wyGOE+dveUoqPYbjWzWZeLohNjO7SnEsBTVyP/WoXAO3kf0q+m5UGIrmWBOO250cOzO
4MG/X7eZ1Qv0H3jNqR37EWdPcChObPunQSWRrwA4XApKgvzJaWg190sB4A/yLP269WBrsEbgjM6R
yK+jv2qLIhTT40ZnlcreNFup2l+U3/szPbV75AlE0UWQFzyD0wnbJagFXDxPH38Kcw3+GfPV4Bd1
uF5fzshQtAtrgiC0rxaVhWkQHBeMTGNgxSpkuhEq48uJsOj+iYjDbp2Vv8rEeaXe4m63m9pcKWLs
V9DCPdG2fBq1yVy4fJFpK6i9xsqBt5d87rdt2VxrGg19epuQGCEXO6ULfQuVGI77vsH9DzbN/YNZ
E5N7uxocr6qHH1nMkJ3+3roccngFmOG53tuos36eDjcgz8G8uAg/v8c5h+QWk/0O26eIdJ2/0GIC
CUah3I4EMUIWSVmdfYW5GPAtDFoFTgH0xrOLXk1s9yPVOtFBT0IUI4Rzw7E2CYV/33V7W1xB9gfB
ECoOdk36uGdk0B7etlwuPEpUyhEMYXBC216CoV6ogbAqV3M56Vdv26rj3m76P1PRq8AsPWGmD27B
fIU10IKPvBNNxWar6NuibaCFNa3gj9QYo/Ionj2lmK5ov+Rhtv186lmUzbXKuqkLNbbTq2Y00gk8
OZTbLLTJufzipCzK/H5SQA0OkfFRwOQNWfSv4S4fx2OieJdj1ivq2WMCtbRILG/IAHWXPir64ASV
2jYW5pOF7yr7sNFzgAJa+6/kjcQ2ssYUrSbuRnHw3qoXj+xN3CkfS5rdCScuolm2fJktYdBpf6Vu
ZHXrygUHOBhvALBE416Rk0mH6fUmj51ntCgl8rhC0spGWJj9ZhMAH5Oj56BAW171ZkDdh2hDZj/y
ZOGMsBWTQJjEOpTjoXOHnGPHOo9/Fw8ve/ffmk73+c/q6aTaCt+5P2SSn8Y+q1ZkjBSlcWtYFA3l
X0tptCgDvotT64nANh/TyTsr/3TyFeQ3OYRs27ThOnV55MNHDSwCSDcFO1oSdqMMO7g0yDQQmsi+
JO9TWE9XdNUO8b0ZuHBP5HFvKExGQLLEOcV0goDxCR2nv/G9rNttf7c8+cUq9HDwK4fLfkAkgsox
0ykpCDNw2SsDswr10HKP8ENMUgj9O0OI6jW2z7RHlSoOwNRAeL4WqSYLS579W3S7DkwSm4vEOmUd
mQUlqw6wyEaE5EvUgroNNEh1F5GFEDpc+5s661gkkJdsWFapectJkO2DFLZlUehVxs4+J/x6ZHmL
nx31QHQsuf410SebfgRGNnbEUH3Y9CMXZANUWOzCr/gygxl6SFx1R5wHNglnHwJpEibkOf63yTm7
5aZR224v2HxJDKQ/CieplgebBdF8EhPPhI2+Sgd6QNQGofftlvoPcFF5Ar/IipljtT85htvUUstE
4T8grVlnkToKaFWFiXGmomXvHWHY3FKqt4n5bUGnE498koDLsY7X0L64eBsZwA3fUXTM92dmPbZq
c1ZIA6sTTdxJ7gCw7F+dcbmKjRmEN+q5ljke4bUVqIDjimEcpH0Gn0HZ3zDnknw8OlD4KwJRDYCH
7fY4iNsGQZIEMXwETFLl02XdvsM/BtWN7rywOQLEEpR/JGWigwJIwB0JpHuZkK7SvvkQkPkQgIS4
JV6vMYba4ddesGpC+WiVebKFP/LeGd6L6XX+jlNpCq7w/9PaKkrxJe2oTnYkZyTjWR6suvyB50z5
fOhK8LTTI6TkPTGyevI/N05AMmG3Uq2utAU4WH2yz5g4+75XMLshPPPpbv04r2aWh5IDNwOHy7hZ
Vb6GBQBq6O4MSNSNOQQRWAf3Tk+S7QyGidDYsokLRDby/Wn7CftOe0jjZmw/nAhZHsYQ4guJvwu7
ebaOrtev8uJxrCJG3gAbATDX6O5+ctNTOGW2662covj6/WBW9cIAWU3j/jUueXORAx43PS9lP16f
O8beq93ETQnmQYZi8Z+Jh1WLFCRajL7Ksso+5cjfR8/y1YCZfUxkBGaaGN7zZw2IZ38Yp/QFk/2L
bD3Gg6+EBTZ/xgDUzhfbBmB+dMfYovxrRDKu/I8PyBEGEYpinXNRG6sZNgr11tC4pCjyoczDHl3q
xfsG0Besj2av/B15Diz73rzOxTUtZ5x/2kZyr28HLspgt8AobGY0yfFYSEndG7CP17T8GWUAMAtN
62/DeZgKhiK/1wqWgiKDqtncmJBJMTaa3h23CrtWgbTOIEY2Cx1JbJjQsMdv9qpww1rib5SIZSgj
7OGAgQsz49eUOuQwqOTWFrVkT1BgqrSho6ZZs50DSIlpFBzHXC54qczY8y6SU8OAkKhWOhfo9lbc
Nqc13MBXd9eAIGMy7Xf/fjdjZTaSBf6+2q5iqPgubogp1ENiHY+86LUP1SClcjGRLWsWd3a3bMfR
bWLt9m2Do+QI2ojG6HL7qPlJiZMNaYjDBOEKzM1aV5rSOdubGgzGwWKKjYH1RMJMs4eGZ1jjW6DS
v2mdR0TlaBaFG5jrhOV2jDkICba4QN4xjzcOhxij6RxDp7XIV0W58PxSAEp4JTubMfOulFHe1YaA
Kj4qCOpPZh+0/ElCUyjpRFV1ZwdOZvEUYEMyD/+wLtqKDeFtlH4xQvbgocxsBcZ2vCmk6fzWa3LQ
fAOSQMBLHD/P5lEJtZPwRjooJmPQMe+Tllsf9lemgXhowZNMpe5n1YhM1KeAb0Yb0TmWTyLAw0ZB
56kmyB3byWRJyoAr4iQ+izcEnfaoEg6n/Z/Xzpf+ofcWF22C61pu4e7nJSPjcSasvUNoAhJjUwvG
/pTnLDgv4qmN93CBUMJSemCaUMI2qNjdqvMyMj8EBm5M2EuQhmKRzj3wqK6qiJhFJ63CEDFIYJk2
eoZkOJl9Zg8OYsIiB1980r9MTD1tis8ohkfqHaAeyr+pWhKIHY0KWgNFEydqjtYOpiMVol0EUe32
+WAgw7PRzPGHI3Gta1mh3VDdLikf+yOId9IwmpgPTWpsRdagXMBqBE/gUTBkyXY4LB0JHfZ1LPkq
c+wTQtaUpzQoxYkHELPPYsHr7e+UrQe6H2hS5Trsdqk3E8YDQfx1Zwug+NaOifiV9yck0THx0qZ0
EbZQItec4XSgTW1rxsDx29DxgjyxyoAh6zY5tFIoTYREOuqxufI0lybMNv6OaW3R1eth+Jvw0soI
gltfrEKkqqv5sqhbcyFelYa3iFq80m373nV7Gha/S3UhVSHOiKzA8giQIJw0CMd7I2+2sdcTAwzT
juIYtyv2FyBzDpXjILO2VImSfNP3a6VSioFFkK4Qr/DlgFp/g+7RWaEzUZpkR52/8gkuA4DiRgqR
VGjFl8NH9x764mHIDhxNGpFlbKssRzI/LcXxV7ebdCcaXaPE4nFltBumedADBvSXjDctCBH6oOc2
CNFEN/6ZWC3dhT3KKeDgokTcL8T4ADLpM25Pnak0rpQrC18w/6Jh3TOCr8gb79WeQyCzyycVvZWo
SNI5ZzOfvHbH/Gc1294wsnxMtkcwAEpjNPXKI1FO16KntmJsXhplsFNB/NeXE1mdmDDEHTFUrQps
fFwZ7xmS4GJuZAtzKmc31FSB82SKVAPVaqpjZCe6lw9dM2+snJhh9d+nYfnDxBsUrQCPX5X6Onox
l3gjxXHhoAQf8ItWgaXAwqVX4WlpIH3iRKPV7T4J76hk52BA7twHet8vyaDdeDNezMpKFmp3ch3w
C8FsdThfTHB/deoZQln4E1ds/PYFMQaglqSJ/ZtNV51QlwAI/w6iwgeIzGfKs+vBP0uaDoGbFadi
DAdN/4tAyRZRTst8O1e1OAlR7gAGjXPwvm2Pot/v/jJVJDxQId8Ncdn4xvGHY/g8OZXDnZetkLSh
fIYpW7FXe7l71z+1abZlhk1FYd1toaEkfYU57gfNcJAXbPgR8d2rcYkSPmeMpi8H3NUSkSP8b1r1
soDsLWz+YMIXAM8rGnpO/Xht4pLJJgw7H5j98uY8YbjLpeOC0WT6CIEl6LYB4mEp2NUBSqzYWpw5
JAHdYg==
`protect end_protected
