��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X��q�{.]VvbC�ޗ�.o>�s��;pp�x�▃�7:��v������)��Kw��'�}]�Sw�����{�* �����>�9=pJ����7�ĚOW���7[%C�.��~*�I.Q�rK�;����L�&���6G��Ԁ4�ف@_7�Ҥ��B 1wA��F�}���q�a9vk���L";V�^R�~C��D� �<����qߺA����xB	�𚱫;��/4.A���{��!e��q��ZHza}������YPZB�u�u��a�nwB��NF^&>"Xإ�zjA����`i���q�����Mh�H��ٗ�o��:���z�KA��z�k� �����*K��Pl/�t��Ku���2s���-W$�t��2�zQ6%����e��R��]-@�_T}�Hq'aQ寽����a'���nUn�<�.%�}��.g�(-�G�b&q�tE�tZ��{�|���N�j�Z�lɅ(�5@�:��h�GF"��Q�7��*�u�e�H���ۨ��ʃ����J�m�퐌������M%nc���4����XW�'�/�`*��Y��΋�_夺�zІe�Ү��[CчИٱյўH� �u�>I�f���u<%�
�AY:v}�'�gO�q���w��8�D�U��Zą_S��tO���X:��Ĝ�H{4ձ��^�+y�V��ۤcaȇ�C"���P饨�|Q���o5���b��/�K�!s�3V(s���E,U�+r�N���>����:$F�x���#U,�5�R�m����6q�X�x���0[��9A���1T�q���m"T.���f�5�k����W�MtN���x�b��x�zY����w"5%�E<����k��VP�^^�t�8/	�r�p�2��7���j�&�zo�]Z�J^��7��J_�;P����(j0e�Rr���5 ��l�%[�ßs �������R�	��Z|������3�`T��v7�8݅�ɽ�A;S�+�:�����zr��)��$ַܸ����y�nW}�q�����sE}u�I㉕��E'���<�P/ )t��P+�!-*��+�J��q�� �x���a�v�0�j���?}�a���`dvZ/�(��7з�
��X�^*�c�tj��dW�R�q�J-|R��C����f��o�跹�ݬUl$�S.��@{fɌ�����_5�N���zG���H����HK��,�a�L[ܵ���W�B8v)MM�
��l;T�
��1����3?p�K�B^7�����]/ҙ(݉$YD����B��|a|��5f%� �ߺm�k)*�~r��&Jn�ͅ���s��:KM�r�����8��s"oj�܄��7mC[�n�H�y}_�D�ߪ*������@;��:�l���J�u7V(� ��'��0����t8���Ra�R�vd���z���vܐ��jo8�(4tU�S�T_��V��!� �C��1�\gS�����;�?6��'�jt� 'e�u�/o� �E�,|�hZ�� q)]U�:L۬�� �c�2�`#����M��0�>_�~�*.�o�v���d�L������Q�'��hv�hq���$w�  ��{q�&dC`T�3��[�]R�7�AH��l��:���y�?�#DdY�	F��i��-4{�&^�%-�]Py=��y�F2�d�C�u{���;A�gI�#�t\|�ѮL_O�=���k���!��8.����Ҽ�δ����P�>��Ⱥd�J�����_�֫C`Ԋ��u�^��O��xk����j%�,�N;�L��@, �ے3kyge��җ1��q�����`C�S��@�u	�'�۲��:#����@���C$�lဪ�`=��������ݰ��pknC�����樹�s᠔��̌���
�Lw]�A�5�"�.+ckv�}��feȵ(���̾�����+ZZ����̡U��[���#�5d
sL�K�+�+�
�ȭE �����A������#��].�F������X���s͠6ZR�=?��T�!���	N��O�B-�O����(C�$�]��lF��u-��g���[+�Ke]o�����_c#[5��AHP>9�C��C��+h"��(,RWAGr��QL-Y�b�{O���3ٓa8Af��L���Se"I[�^�˰S���Iyk_�!)��?�~���~7w5FH�5O~���P_�,i&tr@V����SN	�U�}�����,�ь#AY�+F�$eJ���>��):���]ؒ'�Wس��`	\$��zJ,t�>v��l�R���	R���՘�g+6���m� �h}\��X��]�?�!��R�*�iO�� ��rP��Nh��8�����B7�j9��rL�维v�9Zm��?4�)�g�:<��i�Npy��9/q�=�'��۷����/4c1��T�i�<��0���kؽ����!�H态���$�x'�w�֥ˈOWrk���1�Y�w����X���I�S"庴�U1:)?۞��tRW�k�gV���ѧQ4�O�Ӷ����6�V�+�������.�����00��Y�}�@7�m(�D�.{��]CU�� ?{>�t�>\�ꉳ��d�(�E���<�lQ�\В�W�;�%ah�#J}zA}j��ӄ]��_��m� *ezm�D#e���FzRe�s;#�O��Ĕ����J\@�E0�4 �B"U
�E���-6�"��lX��U�8�q#�t�v*NDD{�poGZ�̟�l˳��m�@u�bލ�����H��Vq��D�'�ș@��f�:b'wY������n\�l��q��2�6��C��D��_ QVGChxR2��7Ɩ{������Ό ��F��àS��*�=�1FQ�/Q��q�m���.Ȯ�Csǿ�� ̃����1T�ޒX֣�6�=&�'�p?� �v����UEUu�k, ��]�T���p͍�6���	]����N�ҽl�LH�%�QB ��0��,�w�/��e�'O����@WMzg����z�W�����x4"U]9�9T�s~X[=5v�-~~U�lC傩C��xTq��`И :v��	��� �k영!Έ�a�6��n$��z�!!x@�!M_;<6`]�m�U/T���K���0�CY�>�n�(�,5|��|w�33Z\�{~8O��򄯓��d����U�\|k��t۱�N`Ah�-V��++�;���"Cz:ȱƍǾ��UL��rqQZ2C����JPc_w��!����g>�0|+e��//7xs�)��l17_��4���I�U�%A���{z(����(��%6�a���j5��܉S:%��9G�9�e�