��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z��;����1~;ó�!E7+ Uߟ �v��M�a�v���]�P9�Hq��;��p3��W�Op8>��N՟�8��i�yM�O6
m���}�r����XD���(�ڠ�\)��:�Ɨ�|��!�ӟ��J�0-ml|�Z�i	`�6�z�w�z�R[A%����)R���Ȟ�@|AOi��1E�ou���A���Qds�N0�MΑb(�pWg�U�D�Gz�E��=�w<K������cxu����X��q.�R�s�:S$H,[�{j9���'P=l�~�AHuj�+���T��Z����sW�n�a�±�O;#pY�����f�I���b�}��Ȯ?YS��d���CXg��ĵ���}�.��Gbޢ-�`�Ta�����}0~����$Q���/Jk�ʫ�ʢ=�����m>U�X:W�,R�����䢃�ǟN֭���(��"�@WY�l?�,���}<�#�I:3�$~z�5g`��]>mD��V�4�9��EԔL�TY�(!oF���{m ���<U&wa�ߊrIԽ<\�� E0N�����]�Ί��
�����JL���c;��I�o�f�,N��A�S�[��H��N� hL|4���[�
�$U��r��˓��n�`#�.k�%=��]�m��34��C��g�x+5f�L��9к%�/�����ͻ����@}~�71虘���P�W�C�7,�9E,������w��^�b�Lq� l������C7�p�+���Ċ�q��7>-z��2(�^�S�,>�سd~��&,���Q�Rxg�%[x��E(�.a�1��cc�7���FF����=���&Q874�ݺ/I9FqYhI�x]�}����ZkX}�e����,<��i;uY��um*�:���Z>P?gh�t2{�z��d��Z����q�U�b�����;��s_+k�a8��QH��	���[L�z��������nH{@D��[*fOo�/I�2E�L�����Q�M����z^C�3��*-��W˽%d�.�l�MN�{���i�A��R�c>ם�PM�c?�E�b����G��ک0(�,��3'}����<W+����qm�gBIDCu�˦�V�e���?M*�����/	t��1 �x���v�#�Q/{�?5��4	����g���/紊�����hkf��"!��'Nx�%�X`�����M���K�5�iZ����.�V�Wz��H}�^\7�6���ձ8jlmC ���apYCAo�l��\�b*��-`~��y���O}�??GXc�8����	��ˠ�0t�y�%(����ːJ�@�Vn�V��gb)0�i�70�p��"k���u}Q1��^�����`�e;� /�]� \o���s���^��:;����ܟ,*�D��̵+�/�l�f���I��k�Fӈ�7D)��g���6j�W�_'O�[z�c�T��"1?.�����")z���atؿ\��.A��w>�֤R���bn��G=�%����7����k%4�d�����(Is],w�h ѧo�=�gQ��a����:����`�A^b�x
U=Z�y�*�é�a��O5p/'W�2�q�'K�j�4��&D���xW� ��k��hg�8��9Mm�<Yxn-D}$O4wW��BN@5��1�3����7�j���@�:�C?��W��x�4�A���;_:�i����i߉��v�(�ԒRK�����[rT��x�/g,�MJ�[�/&����v:T�N�o�����gwE3�C��&�S����8��=�T�j�ydK��H?<���2a��O5 �"�c�@Y����@V2��w��pO��ۭ���Z̏�]	��w[�q�/��P}�fa%�4�WV;|����w-����IvT�������x�����$��Iz7����P�WH/�G�J�2f�zM<_pK�3���.�6;}�&���~X^�"�P��^�aĆh��
�W�bH�t"�s���=��j��ۿ1��Uٯ��O!���3��XKd&��{^��zT=�;B���G��Ur�V�P�-���Q�u�}��aK9K4[1�0��@��f��8Φ�(d�ZGu)��r�-�>7� (����mE�NL��0GO���
�s��RR ��һ
��"�͹;E&�^ސ�F�Eα�E!�p�t����*�#Nh<�8VgZI���[��]q32 �Ҹ��� #�hʜV-hn"?�Dd�A�/¿z[
N��"�$;|��1���SN�AE#g(��&Ļk�1��F��{�	(��:]��{8ov�b�K���v�O6���t�uv���6'��վ�c��F���ˇ989� 7�k�P�6c>��p��I¶�u��7���fc�ˈ�ϬS�@�^2^��:�xt&莦�J:'�g�����ᆂNcZ���������5��@�%��h�$;з�9[>�p4�ǫ���7�WY�
���:U�D�򒫃.�w`@g~���L8���� �â;�թM|@|�	�.0mW���n�>x��ζ�KJO3p�a(Z�ƾ�\�*��F;G��WRH�#����������Ó}֩)��� ������ۿ�_
�`hB�_��n�,�[��x+�z@'ɣ�L�t.5q܄2(xi��td�!�D|+΍�o{�z���z|Z*gx��?L��zz�}{��U0�������O"��2$������UH�_mSD�ƊN9��1�#��R�.�r�&�(k"Jߡ�^x6�W�e!}8>i�ӧ)���������E� �d��b�.'>uyT;�d9d���z"j�]q�9>�������γ%P2�/$�����T��,��WxN��!��/���F��Hj�OSo�D$�vgDAt@���;P�;��>�5�����Ґ�	��U_�̅�c���9���2+r�Dܣo �6���[��}�DϘ
^)ؓ��ϴ#=u2��*�R���?n�X_UD���P�V�.�G��C:��Ot�	��|�2<�����hU��*e�=�⿢�5�g��H@�B<��y�v�U�zj�W�7�tP�_F���9Y�z�yLK��]Y!M��Q���T��=��Z��_���Ϊ�H��%{
n��@�Sv���!Ɉ�	�H��Y8���@ߗ6�B���su�5C�b�����J���oy%���q=���B�*nW&��@�Om�1?�M��+3q�V���|���Úx�~�Iv�������vَ�k�ΐ���6Wۭ`�$[�O}|*�R���<̂�ؑ�ž!r���� K��z�畈�嫆z;Ǟ0�I*n�2�ݤ��u�h���g#�um*FiR8����3��V.��>��z����!�ڀ=m���C��g��;���Eo����M� Ȑ��c:�w?Luz�EoC��dS[�o�g�ba��:��]�����:����܇��|��vhCL�$�#p���1��"w�%�شupE�����o�2r`) ���OI~���:nb�.uL)���,�.�8Y���u�Ê���'��Y��:�G)����=��?/P^Z�*�r��6p�L���@{K�ʂ�;�oI��"���ŧ�@�P���� o�O7C�"��i�X��b��)�拭8���_�`ҿz���/{�&T�J���⧷��������K�Uo�I��˿�<��^�a���c8�gN_�cY�u�_��c�S���껧����6Gw~���ͷd@�m>'D/#�-�H��G��a]�G�1EM����[� �y׼i��xg�3ߪ� ٯ8��ء�+�m�gÚ8b�.n��W�����xm21N�u�8Zg�`ƧZ�$��im�/�o=���$�o��Egy��-X�}�5�O�9?8�H>�զ�P�sz�ݚ<AaOM;��}��h��4��bq���ɬ�aQJ��\He�)�M�)���0�H7��'��k�ö����f��Mt0�C=b|O+(�ǘ9�Wn?�T�O�L ���M�ꜧ�g�8 ��N*�5�|�}�DA.��t�����,�*|2Rknh�Z}LT��Z�W�������k�?	E�,��,H��!�O.�Kw�3 PPJ5���i����Š�<ߧj��w���g̠�]�x��!O�Sb|Bbj�ݻ��5'��E0I�.���+&vx~���}tY���5�*���^�oa�\��NHn�uCժ�ڔ�d��	k�m��R�����1WY�Vz��;z���Fc�ME��,WYD�	4�����-u��5����տ|�؄���x�򺍘�X�+���7�F�NO��E�[�N�ZaZ����E���� �����^,�y+���{��U 9��v�wP ��f���!Y�ʴ�JC�L�V�������d��{��-�}�yJk�W��,�t"	���E[�*��@��osbB��Vm�vK�~��哜��Y�.Jq��T��A�Y^�Y<���q��$� _��2���e��,��=6�-U�X�?6te��D�ǹQ�����s>���jn(Im�n�[}��_C�  ��.𭵟�G�����Μ�isy�Qn��R�{���,���0Ze>6Z�F�X�X�c8@�&uw�jM�;�O��S����(&D
X��t�������L��r���M�1�'���J��6���"��M;�ׂM�Z�fs/�s�(�Bfe�j�	B�j������Z�O�B�^˳@����h����*�����ҟ+��fK��x��H��{���J3B�>,xE���l�A�[ɻN���C#��P��<m���<<��P
��܅+�].�{vHB�H���ϰ�9~7�2+��)\��vH��Y�M0�Un.&=F�6�y�4fm���Q$�-�6k�x�!�4���V��$�f�פ�m^���?�kM@7���\u��6�a��qB��$�:	�O�p:7�rp`"�K�9j�R��]�7�87L)����C8��e��\O�Y�1VV{=�6���K��P����1��?\��'��D���B�.�RƜ�w���K�X0kn捆،tA��m�3�X�k�y�f+b����t��)e���C�ar�މ����"�y\()-�M����_z�2`����O��L��:㭹��'���J�V�0���{N��#ʭ�f�J/cd�/��y��w�ѱ���?u��2������u��e�WȊ���6lr�e��Ǉ,��Eq��5��C%����͏����8�b/�rt�v'H�ل����/�O�=��|��/h�CI�K̎iM������c����)N�#-���[Y�.w�cҽkj]O�*��;���Y}�čL�?=��Ƅ���RT*_�ED�!�ZoSzn�	�<��}�%�ěL�-e�V �."�-Gh��g/y�Xz����p�5|����'�3%Z�O}m/a����dj1�m|➜*,�QJӼc�,�J&���8�H9�G�fC�����0��������e�T��w���:nE���`(�B�m^җk��&V�*˾.l�C3J%\U�6����\� "/r@}F~�!��Zht�W���C�w	��O�c���ܬu՘w-@�/�M}���<d���qL��Ԛo�^�L�=�PcZ�Ma� ���S(�2M?�'� ^u�x�4�oq�,��h�J��@Ҍ�۫-|jm�"�L���)"������FDGE�K����0�Ͻ�^��lR�~mX��[)��������j݁n�t#�8�$U��!u-�Qp	��1 ���1&�-2J?�����`�*����5s����Z���?�NLd�HO/�W'Ʉ�L�6eDLq��Ha�Z��r'3_G�ݚ��H���nZ��HX#`�	��jw'�0�rI/u���P��ۡn�ǥ�LS�zhT��'��ݱ<ke��\�iz�
t�/��=@���$<�8���܇�:��2k�,`�J�.��g^�"Cҗu���;A�{�W� A힁<�yXd���۶p_K0ފq��`��Ѡ�*�!�b5*���@�N�]L�ѓ��{x�m!�����H�D3�ύ9Sg
f��|% j�'X�1��H����[Ԍ6.p�$�xV֧���i�=i|���ϝ"���`�i���&�}���Nd畭���K#�>�o��,��r�f�wqҿ̴8�v.x���$�[f�J~u�XU�u7ziM���|a&�d�3�A��[(Mʡm���W����~iA���@Ī�AК�X�cfP�u� ��N)m
ق�_�[y�*���.�@����f��
�+|7�^m�\�7��ݘŷ+�
y��9[EwJÑ�KM����U�)������gk���ә�<���"��@�혍j/�5L��K���<0�� JĭX�� +�	�s��h�J�?lp��t~�Ǫ�Wc{͉ �y�
m�
��9�}��EH�!�V��8.d�����!��n�k_��,���ð%����Qb	��ɭ���N���4B*��i�5;J�O�,�����5%{��w=�D<v�*����sj J��_��'�{v�G��<���Ry�N̐���z`�\nbD�`��G�^2�q�l6RZ�p�)�;m����g�sA���vɇ���.
�o�q�'�օ��t(�;�p]-a���@��ި�����m5��slı�m=��Y4=@v�?���q�ʅ�2L�%�ڸMcT�&��ri��15�����Ų�c���g[rQG)�=�2H�t��� <�䍣7����Z��Iߒ!x]�ኰ&/�t�ȯ�3>��~�'�d$HdDa��4*��s�5�!γլ���g~6��\DS�	~v�KKA���aq���k��!�Q�N����S�����(X�7����t�]��)*�A�!__��?�R�n�R��^����n"\c�DZ���Ң�lh#�#�(%�j����fÜ����+ȕ��������y$3G%��٤l��?�~�6R֦}���5\��)���z"��^��͸�s�>T'6)~��"0O�	�r�����T՟�?G.כ�)�2�-F�-2o~�(�>�{y��֎���d��"d{ެ�f��S�i|r0�gX[��V�#r�(娺�	R���[~�p�^GU�-�0e���S�������� � %����U�=����eY�m��Ə8����Ue|G�ǿ�ݫLq�d:���a�П��S��0����.Ρ!�	UB�4z���?�aC��Ƣ��<�c�	����qD�`L:r������R��O�Q�8�`{k E�3j�-�cԈH^��3 Tp�A�FC.-��p��ݸW�O�W�,z��X�,��vug��yU���~2g�O��(�PD�z��_�s������ES�!�ͯz0�I��=��
]#�W7/��f��Ym��4�!j8ep���LF*<w.�VI?�U�mAtn��˕7HoZ�m��s[�b)��Z��񴓬��8��"�#J�t��H IN-�����%�\�ޮ��Z�`{M�&�|S�֩�s�Y*	�QeWĈ{�aˍ5W�����o~0kDb�fK�	5���k�Pw���k��[v����cp�&�.�R��`�H�[ñW�H���d��$
l�sa��\�]�x��C(�G�u����+���.Uww�54o��5o�.ITIGng(�c���ƵN�Q�@��6���.�k���%y��'���K��2Q��(G(I�������ku�d��3,���0/`o�����d��>�p0��3NM�@g�`C�X$_f-O�9�0oL�
�3<��*!�o�	D���5vs�5<N����/�/0 ]j�]V�L��(ؽ����O��O����H<��v�{<~}�%�0�Վ��k�L%��H�M�_���#!)�t~��w�>N�V��ڏP���":f�Ilׄ+.�Ò_���V���z�֜S��!�W�K^�Z�3���{��
��}::�U]��9�q9To����F,�}���Z�,:dc������������@���96c,�X�+0;0?9<�2��*T}���~^M}�V���l�Rc�Ϗ���C����� �(��`�j`́DuF��I 
!��h��o��q�8l�����4��^螃 G9���H2�4y�����`ix�� ���LP��\�u�(��d����GrL֓V�
5!�L~
?k .5��z��ϕT�W�~`��:�Ca�N ~��E����BF
@��M�8��#�Z���F���n�Hn��6�YP��+X!d^�^��u 'p�m��%"����?$2${����GvV�{�t�h��^�^k�Jn)�x��MHk�3�,�a"q3��թ:h�@��_�C
������;�:�n�p�#�{bɭ�Zs�P2�ŔGo5u���z�L$ ����Q��@�&�b#R��n�?>o}�>�b�:��,��~L��<!����,�ks���dI�N��a��T�%º1��9�Iꗍו�����-���!$�Km�{�p�� �Sf/TrD�0�Ġx�����Ĩ���P��L~�����yG��l�x��%�jB��'�An=�R�\s���� v�K�'�U� �G�����U�5�z>��сi�بy�W0�+�s��P&t����6?��$����x���3	4v�>ދ/ɢ1��C�n�FY�������x��.��	w+���n?ц��ďV�ɩ���|{���۳���rJ.�3Y�-��I���>۰ez}G�z�;��?����kT����ܱÈ[j�2���r��Ud��CH+���8i��K	�w�\Qi��7͋!�"=HC��)�*0�v������A=�L
N�_���W*�3ڪ�*����mc"���71ފ�dk5y`�<��B��X,��}��W�_��ѱ�z]��ry��?&�(MB��"����q��$>�2��tC	�/d���0���e9>^T+�m��Q�l�|���#i�	)�1ު�+��F0ޡ��۲�X��3��ue`%R��Ѻ_x�[�
��jA^c�i0��d;���$oe���)���������/�e䰲��\BB��z��@�Bb
pqG�f�D�_��>���3o�@�Cc�$քy�d�]�C�Z[Єr��:�'w���0AG��I��a�0��.G�R(�QsI@�?d�у���r@���m�Y�lb}v/�cpm|�'�E�P���OK�-�r��PٲYi��mHQu��/R��d��0^��u�vXmb��ߋ0Aq�I�g��3�b��ɷ:D>��[����V������
P��7�BS�Or�����_;��WןRMo����`:*q����|z��+�ۭ���/�"I�،^_'ګb%@���#/�O'�x͑g�����)���]<�Pʑs�C-!��c
GJ�Zŭ�P��@ ���]�_%(�x����+�(�K?��X��]�B��"2O�=[+�(r�ؒ�`F���6K��N@���P���\5�7�(X�֢>+CE�?xq�kf}�yb���`Hϋ[=��rv(V:�ҭU��7o;���.� ��}�k�u�$(=��2�&)KֹԈڞ�Ʒ	�;����Ƅ�s��e8��7���L���U�CC�{�튨�(%����u�M/�q�2U56jJN�1kSS�f�6��[2�w��lb�f\8�*��_˛�~G�	�Ěw+�+H"��Bl|!��BW~��g
�`9{�Ct�)�#S!��؀&!��s@�E��������CP�����A��n�V50�Bp/WMcW���	)v2�y���ܻmP�6�b��{5�����Շ��n���[
�U�H_�2�
e�΀�UZ�$킍���|�-��O��0��`��N�n��.��D?�F��������nMٗƇ\F�Bj�^��[d�}V��n���y*)�	7�>��:f��׬�y_  �[l$�ksEj���Y*a�-�R>�1��:zါk_^p���#�C]�/bO��Ub�*��/��Ծ�7���%�;;��{7�@Yl�N28�.�&�i$:p��\�g:�>�<�'�b�I{8�Pb���M9�ɦ���ЎR���uh�4���;����ة��Խw3kt,;A�W!�W�R~�l%�Pb�-���)��'��-�(7�x����/�Lc�_�t�{ �u�8��1d�v���nL�:I��C�<$�����jKU�;T�hLD��x1#�qxI��h'���-ⴥK����r��&��Y�P3ky~�LJޘ�k!��c|���z��s三@�͙7�M0�Zn�~"��٘,����-�p��ߙ*װ �6J"HH���7��˪ݟ�t��L���`$�,\�Do��������y��yH��6�8�p��A΄���E*�.�_�-1x��m{�oO����v��L<���B��N廐$�ʝ��"���;�,�v3�J�p�>{F)�2�j8�=;��3�a+=̎��ť
_H�xr���sFW��`����r��-���6�kj����%x��������?�\�tb�2;�3s��V��A��{XГ:���]�$0�q�6�S�ls���]���YA~�I����2��4J��Z���^�[\��*HY���;���?3AP���1��iy���;�rE����Q�?�xo;�#��(v�{�U�89V�`݁<�O4�C|�M��t� [PC="�'�p� ��(�%čv���~٥5�����K� ~�v�����k�3��8(^���Rl�C���	[��� {6�/���B@�t�ͧ�[�Ũ��)��8��w7�1��IY`pBs�h�>����v'�ܩp�=���������̭}X�u�p "������c1�R)Z_�ĩT�'�K�|}߯J��R�����-X;' ��\Õ�x���%tE�|}5ř�dz�
�a��RFm�Z����t`&����V9���%�3����[�*���Y7���c3�i�#����\ 8UD&GA��,s+c��*����b��A��_8K
������rL�s[ ��KYjR�X��Bڃ��8��id%pf�2�o�q��5O�
�n`5Z�aa5�)��ʽ&^H�)�
�e(?U�j����O��0�>�0�����pv�U��P
���iH�����K����>��H��
Y�d�3E���b��/᧽����30�p�De�wk��0��D��kJ5f�(:KӸ%L�KAZ�kiah�����9�I�F��@B�</l��J�k�\��[K7��?�w#�.gu�:>0�)�܁Y#l��Hm%t��3��D�p������F������ ��ԟYB��
 j�!�D�Vz�ރ�r����0n���m5U���l�%�����X^�G[�fxZ��0=$��B%��ܒ��ۮ��J�/���9���=b��X���cVi���_��Y(�O� IDH␹:pW��9d�����0q��q�K�. ��m�R�MX�����o��]�5�j�6b��H��Ʀ�8=2h����]��<!F$�5H��@c�8YV��?�ڠˋ7�6�) A�۾!H%"�ٝ���]���yT�NL{Ϥ�=Pr��Ƹd}o�&�Mz�K �H�0BD@�_��1��ӿ�@�aHOJ5�Oغ �K��4[aRx_σ��=֝�v�Қi�P�3O�׌p������W3ˈE-I��^W����·/_�)�Y��!����γ��{��`�"E��1%�u���9떖[	|��l��W/cS�ϫ{
��;�@��Γ���E-�����%�����;�֜R�YHc2�wlmտM��l{ �lÞ�L�/�+�C�{?ށ�dگl�i�	ξ}���gη�� i1�|�1����PloR�*�V$	�k�O2ڍ�Ë\���p2�~B;ѵ����J0S6a"��]�]�ڊ�$[<vr�y��cG[�?$:�9E�W[� ƽU��-�ϥ��ӏ�Ph3�L�R��:I��mԷm,�7S�Bʔ�0��CA��:W�f����M��ASv6d���T�JU��׃�2�B������s0E8�� ��i9