-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fg2KcU2DkTF7xAmUSgZXoG4BMGAZpbphBwQD/yZy52rcvD/Jz9lYfG1QfAprztauZRoqA2izE2up
S97PWGPO0rw9NV+O9kSnaSKLiOgAry+i997+woloo21qT2qazdY8m57Cug/YqHQFsmnTahzeXLUr
llxjvxD/suHQD2+9u6SrzwXEgsMaP9Swi2TPErNeMa/BynQXdIKmdFnTj6p/socm0Z/9XY/fu/ZW
aXENG79/8FkCo7jBHDPauz1bOVpl/UekvJjEltOV07SSUlBGP5BZ8lDfmF7spfUoUL/GBCqKzzkg
eHvIUsfX2TD9Mz2r0WQ2/p61N9K/A6HzeuTy6w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
1Kwye2aJ1EWZTixWVukpfqiIQkUE6HbTdIDRKZy7ECB3seIWOh+XStlwV+H+SKbeCyEc2MzgplDP
Krvu6MnY3AMjDjmjzAK1cqyAq4p4AvZ/wNN0p/Le+j5EVxJ6zFhixkiX7xmE4te46Uo7y84YAqVZ
ZjBdub3+6WgbarYkIkSU+WkwpCr72ljUT+hoeAKn1Lb2l4xmaLIzwakohCpBFedtEaTiCoqD1lbE
LZisAL912xW1nIr5W5feUdO4Xid1oUQfJLqiRuGbnSAn5fVDh2s0bG6IkTHIm77kq9NLz9irE5AE
KcjPpf2/stoFyHQCSx3Rua6q5oUs1pBxoe1Tx6YcUmMckIOMRUioR+KLsuujvSFLPoMXNcXZbPaF
U0YVhyCyGhdlX7KJTLOBqpydECPoRnOdqaa85/awRBnFP6ySOK+RXHb/Pnmg9lIDye19RozATx+c
cJ6VKeDTKNAvcGk+sP7sxoV7KxKUviwaXIcFCk28KKG8lVZ6pbF2652+fQnZ/FUiz1rwa2q10bSv
//mZtbTq1aOhHOSO4IjoQlDdq+U1/vsdMOKOmwlfmmanVzXkyzafHKclELMe4ujKk77UqwGP4lgP
c6bUwkR4d+ola3E4Igc3Kghgl9+9FGh4JeDrVsAykUx1em2CfYB0Uk1En7e0YsEhCS/fdp5BtUT6
6M1wkUZ1zcceO38VmtM/1N35Cu/ACPLAF3OtfF28ocS6ccLqMAOEmXZA87m+655c0gwIPqMUlkE9
Qbf6GMasj1RpH/MfsTBdfKwaGo5KJnLbbDdEXDvZ+fYyu+eKv6dHgBDQK92zYYryrQYJkCv5K9hY
WZ5mMOai+IVKlFg0Ta2XrJvjhvzvBT1rLUKeuCVsbtejoTxgpRKNQFXZxsLwLQeJw5/K7UxMm/0G
Z8T4c4hnOEz0UtscRNXoCQbXJZjD5UkD3I08Bec/Jf4/xgWtUVp3uAPudP2+cdTajCmB66z1p+vG
45u0bW19OtIxLoe+ugp1hUa81d9mr7Jh9VMdAjCxK1J10U6dLQoluy9rh9vm2iFDP6u4gnHzb+at
8DdR1+4GQzGC6qEQ/9/mVlAWogqgaNf4pgOcAnSD+RHLa0lTQVn1BU1sNvxGGFwbxCHqiwlf2WTm
ewN3AhnnD9FqmTSCDHOusVoGZN9ucBmB6aQZibIkTs7juUdPUIHx/SuM3PD0E37oexKD3Yj1O/AE
NSSXy9pbEvUJkdOVIudb0FDtZ9KyWxM05a5RCKNt2OpzGv0rRTpsZBrlI/xfMluEKPN5SOj72yCz
iLWfA6BvwP2gxiRisgF+HsblhuYqw2nXFji0jlHelzgMi9GF7415FmckJ9F+/A+46rtTWRG+UoDg
Sy9tuwcHxwQXvZh9Rvrrit4LlWZ3xrtpe1QPBDrDkJXbFsOYpPpT/LcFUI7wzckgX5csMk3ygCKS
53gqFiurRFl9cTxAqJs1Kawriosu86iV0nGDAW1N5p2Dl38XBBcAbu9BY5sTPHSO/QlPk+hkZok1
y+y6To8kcsL8IkNQwQJDxXIH/j5ouvow111TBdoieOHka+p0SboErmzRGz7cI4WsxSjINeBDizxa
A3hZDo81/mw/1jwrWObHr9hddx6ycGRC7nd2hBC8N9s6te7xUflBu9l5uCkz7w2Gn1FFxf2GqKlJ
/AWa1SuPIYUZA72zRIoCs2pZ/gUrNpJyF8XNfXh5cHIoc1YHMKK4w6c6LSrnFZrF3DB8VckkO8f8
PoZWxkJ01XHc6OFQ6YNQftKwTY9ErbKzg2fu3XhRwWI1QcVPN1hNT5ZZQoGGEtNdIeCmgc98qZPm
ZupO4zVldM5s+3vImrLGcSIIgUm6X0sPk3mPvUNz7eCSX52SGp2R4oZ1NDtB+Yc0MXCDlsazgdBx
OMpfBd2Zgp+6FBDZBsuGQfTJMrSb3XEjbFku9qht5MjvnwA9QF9GtMuM4RMsb3yKZajGE2OKtnh4
rZCH0SdgXfkrcI/+Ccmg5CRjkhQBJkgSFYz5ZMkIIOYi2jJzKq3Pi1VUAeozqbOHKsqrZWp0znIU
OSDoV67f1Wtj6YCyfVw+2NG4DZSJ6Z2a0zR7CpN6+mGRq587vLOSoO/LDTM4slyzE1caeRb1CcU3
whH7kwoOIbgb9bRyXOQ5M3MXXD59LfArK6gFfDGY56tXlrB/cixeBH868IvAoEGbh7vgVl6YQs3V
naQqknoIFIiyK88V7F2aBadBJMAYu6vpJeqIBH8jxtijc3813fghE3RldH/ROBMV2d/YJyLCQet2
nZoggxTHwCi16JVCxdhzjFPr6h1YF2G6cV+OHImuA76jyYGxVTGbwWT/9iU9DpYFrsJeIli39HeZ
9sEsrrefs4aeHXlKzdMIsfK2+3zztBeteQgjL915Ycxry8XUrOj4TyRGVNV2Ae0ciAx0RLr9br9w
F0AH3dZ4+y0+7MoojkxUdXm4vfHUKQWM4F4wUrgLcxDIdK03uLvr4SJjM/f4d+B0Cvq4eXFSgRkV
0vd0oyvxw3Ecm+DbpJj+pVUUx8lu048Rwt2pmiOd1/fi/0rIjQhwOVbwBD7zJpPDYVR2qsRYoF17
RWd2UCLuMcciUqkEwtV+z/980KWCbE8BoluCeoEkzyGyYwU8h2tSpXPj3TcvCrXSow8FCQQtIwl9
/h5O6DoCIfUmxkB7hdND9gqDJW3bdoa8RqNQ/pjk2KA891gLSt918YuQX831zI/wkoYfcb6heYeA
ZYFroDzhLCugziiBNwg+wrHiFSy6IL9Fj53Ta2jnYNlakkYfuNL58DYExPZPnNpUO/V7oKS590hX
0eUZ6O62NByntXb7r8ioZU1bHl5/z4SQWssP/sIVUFErihq7XNiH85TQ9eLlTfCHwjrT9Jn4KkOW
9itvv/yiWm3XwNibFLLP/n9znRfU7zLBzDbIRK4nXj53ZWk1g+gLkYetwSqLHd/XY3opEUu6sI5D
t7k8X6e10Dvo2+vKUYstk3PphUkSS7UhaWb4vpDqzRA6m9cT4uPOfsELZ0F4Uy21Eqw56sJvdHJx
oQXH2OcU2zx5uKOVeEJlxayFTL5gECbjTI3h7pW3mg656WCKAvqUG2kEi+Jx+22+y3iwjMWlM3C8
kZ5GGtbwvbSHym2zdOvJC+hyAS3z8Gt/veg1UzqaUEmhzQaUamQgKrDNMUO6B9GIxxHMmESht5oJ
z+yDeMztOTUj0WhmxioT+hf8pMfCU6/0S8czgaV8RfmrjcN7fncRQj9/5OlKqMp3Rm/2n8HccLG4
fObXWyOjQ2L0zA+TqZ9X5z+wJN0fZNTL5CFkDpf9g6HWWYwcd/x93EXQbfsBvPPUMvzNk0f5V5nT
S/LrN1FLsF/dsNSZcihK30dBTucQEEWLO8+cF2UmG9YeqIZUF2jyL5FFlMloW5TbArWWSQHIZ+aP
n4rxxUM8vFjml9p2nl0kEcV0xFYP/fj/OmlMj525DlCokbs6gTTfuVELZbyYO00F8wwQ5MmMrFNP
YorM4nxRAxwY4d/5BkUuIZQVHjKTiakzi66JAG5sHxHyBki/6r6evi+J3H3eYAc764UWLFnCsL4K
FeK84p+x1c152DX+3NveCwqFfJHRGs5zQoHTxPF76MKBhDTEFAQdHfUdc2Ty4rsfqIk6/vL7HaEK
irdW8GZjabn8QQPlw+mrzynQAw6DFo7FO8VlmRH7vpZcG9zHdxf7AfcjS6l+7uqG01nLRx6GdDBP
KYW/nQ7BOv5K0rh2mIXj2UJ9sKZXpTcRuBvKuQ1e8Q8VE1N7sf1vFnYY7jMzKkPyhXFy7eklegNq
9TFFxl1fZXlZToSWemG73uRT7zKtXiXg/zjJ64p+q22ZRJAP05GGLUtv1W//jf3b81PwfuyiYLb7
bPycq9HiMTd6D2ARE0j3pyXDttY9zivBa9Cc8YW0Cn7DyxxJTTPwYtaySnvmDRhNs0iO8m5/Nm16
Y1+34ODeOFY85Ft6SMrSs9I8goNQNjsrzbRp0aKjdU+W2+zGuWcq/g86Q1r+l1G6oNVp5axlFet0
SuEaxn/3ATyNqfS+zi81TujfhnBEosls/lQueFv9I1e6RCc5sDhIeHZQYWuLbLdnBtSAlHt0cWjN
e43xtr3+WlM82ooldJBzpnpc5iUk6T1xuoLOj5jxZF4oUc2hJcBIfYuglJ0fYR1ltHLJGYS44l4x
Ruf1TvoHLAScJmuIJi5FoaN9wQIE0th5bM5Ezz6wkrGt14ItOgANqdCsOLhkBoFfRJ/9BG+U72VF
2e54iQBL1CBXS8e9hh6YlMbAIqlekM8EcWl7xwmuTRUyLmphvuOK+cmula4MpVh8j1s7aDJD7Y3m
p87kMOjvZ2SEdb++0FTpjdO77pB6s03nAuu6clTyxfIdooa4q8EDn41+vKOn5D/ytMLA6gSjW8jP
DITVDwPFWfOkx4C3BRZKfTaaR5NOERh14JEF6tTNmODRhYAMAZKV/iGC3wIemKFbL81Huiay7L2l
B5W1hIuv9wJetEz2jAEPvT6XROq+ueBJ53IILqMGYmLiCMbTwHa8XuTl8KWmsUKiizuQAEUdUSyS
CXW60NDrwrMCqOKwEhj3rgpl+hJ1WvuAjPEdIpMixmYKmylr3EmWFMrp1loI+ttXEt4rJ/3PNiYi
l/LnwZjKtL6oBEG6t2ZlTX22HE2BckblFN5Tn14xf4LP2Dg7zI5/x3OL0KAMAx1LGJDdDDA8KGMX
LcCaOcnzro2phigbXAdWZ9HzGgY8e8ESjYfgVmaCSM0eD0jjcFS5LetNjIFxJ03nJn8xwbdpzfqh
+VJBAAEe62ALzcvgThXjNL5GbCWypBa1HBzvgVrQnEuS1ZQ25M7fJkNNHWUTcjoXLgEQpVtL3Xhy
dnrzJJGkvVjrQZwREIqY15KQHA45PxZmthnFakxYdiJBb0UN/v6qK9zgIVzmciy0U+O7p0rXTo/Y
y3Mu+rH/j1hF/ddwqbebmDQoBlhj5JddOWKyGdw56XMsseCbPL0PoZurKbA9c2s13ldJVTe4R1PG
IBfWhhzHnPIhMoUJ8pCGUd/R7eeEAGYsHkl+Zy2LFwbvBdbkzGhomEP8A/IeHxvgORplC7JO2cX0
izkP/XtMslWUJnWZG3rQ7+KjLqNB1B0uHIkLM2+bL+ouEUjtvL00Ep22F0EJDFgMGjXAcHMsa2Hx
DMKblA3NLtvWKgeYzUysvtJ6K8b4RHGdjESrUOiRNLEAiPp7a9pkxoRpw1A1SpEjIx4AvNsL6EPr
uXlLTSXqC3YE6dsVJxrFDLqhZzXdg+4Ssh0tXgJ2phO3ASisDb9jybhO+Cqq8Te0D6o8GD2ZoXIY
cehcNuSjOnN6083PBAH0IREPqhk3fUiSIzMI4nytF8g8IwKAh4ituH4EDuUjwLVhpEif+Q7ZIUk9
5Za+JBIGyLrDJqjWyLisARnsLP2XNKOQGaoKrQDGur03pHHLOYnKIHZN6tJ5zf6u2C1VVAplQd3P
bi7jFRO+VRNlB5D9H2vxAar2iRFPF1BRDF0PAADMMdsNr5O56id32xZyfftsMIq+gPgzTSGWeWjj
ccartbvrg3VVtq9THlXpXcyqCkuv0QBTlli/A2bgCgi22+vV+77oPIgkotKYdwK0owCM6QPRiXMX
2Tc9n8L+adrmpVAnehNaWOeGWcUTa48MuJE5SccLNTw3Ebo4JkXZE8kOP0cZVu72bt7jzmaKtkv1
DzJzEPFjTsee7V8sy3zf6PWUU7geC6+gW8vnD0ALgF2sfqvChbGLxqur0kS48/jDWJxUTP5voen2
sKeahUDXtQqtgPvtRrEDXClhpW189EGhAOx5KnBMpTAcvFKSNaruWh7qMdl64PlBB/3omszMjPiu
hZYT0PJhbh7jBMo1IkLljUZA/YaByOBvwP36tPkXQVvnvz058RUpA77VfJQvGFdr8JrVhbFkmqnW
3h0Yf6BkFVMHEhXcHrptbuWPtmSfS3v6ubFMuwupEE/9GMo8PMNw8A08g+0hMnZlmnhexz5o2hus
NejlDabXZwEanu7IH0QmR64DkNG3rxY3nQjjHX8Im0KvKwAe8+Eq7vlGqlm59cH7e8dqxG2z0+yF
1HL7UP716abvGT1Zf5EIxhOJ3vmcRi5syL2Lrr2MLWulwsbHV8GqjyqjFtFWEK6fJaxeH1FD98iN
gxHN8J0kKzfISIpM7qMhnYwiQYYgqqpPmXDTCeaXA10EjhrgkLD8G54oi1seGY9qSwCPZScQETiO
40MaGalMmvibDhrTTRpqoIlKuCrWeXz8vOrWzSbyZSvKJ6fJcw6BJ7dCtTGxPhbmy8aCjb3PhfME
ErlZI2yUw9sieWAUlx+7Z8h2x5VA4h09WByZpBpO2qRJB/RFHeoaE5LQN2hhMyDwns1ZpxI81+MN
xqMlAAqF4LachS363C/dUdnvHYQqHV+D+ppFriqbti+PwedEMAC9Eq4IBPxDNLaJa53D0A4Y/O8v
Mw9l7jsJOj8kWMJNrb16OXVz4tT5Uyf7aoZB0HZluSeji1dkF+P7gknAEuUdDgpJHiSe448CNAoY
f8niGwEe6zmSRzLo77qkAJaYURGCrAP1KXiGTwLWd0ryWVIAWzMpoLLRNPa/4yIHzsFIaW2d01yX
hzXVoyNC7idJ3eT/usDr/8y31lcneAQ5CmRVxtKpWJt7sECww4hzXIFgFqfW6djtGJbrpfPB6Ljr
wor/NhZAEGWmExRI1h1O+aWKyNfKlGlYVoa+Aaj51toM98PkMeUfI0m7zaE5RkEqCVVshRIVorgm
a7OFzOee6+wDMAxrEExQongAqroJ8+iexNzJtqjgaSEqiuTsFRvrYe2lXNcW5jCDoBBb7h6tMM5S
7MaAcjm6NRMkTu/FgbHGGzeskxJSLtSy94PT28vvKU610Z/1oAkE47/oetkfHoEYStFnHByJdL5v
bFpKJTcaP/ctwWqbMinnk2hiH/1w/FqnGomr4AIrFt5RHAVJMsjXRuvg4yhrWR9z0dALyruHDGwb
/GgEgEBgePFHpcVaL66cpQdG8qvayTBNxrDmBhL6DJOAIVPMNTM+3IxodHMaxm8o76nO4WlPjA75
5d/a4DWpz/ymbn6CUokCxyjm48Fhsu3A1YhEQzHwgoSR/PzENtelTAkgm4Ev3YyTNgafNv9lVcni
/rmg09vxbJ31fvqWA2oTVW+OUM9oSpZZjHmcIhi59sQW1KT9FHSQ64txSvxQg1YjlO6r2NhYfSlq
lI6sL2+OLDkaJF+4KkI3e6NoUsNlMzi00ahfof0xFEXGpx3HAoH8wfBeh+8PxO5nfji8xnhoDX5H
cWuE/kPB6sef+IZYdZzwnPEd4gDCSdTPky/dIC5Cky1E9ehUIOeKhu5qVHYuc6J1wfgk4cmYvDXD
TdnIMggcsBrzVBxMoDnoJTPAxo19eilQrbq9Yo/EQd8ZfEu3sfJJbdeNFSqGMMFWPKdBy0Qop8Df
JJqaJCz1lL7YtuFrDoUiXmt6h/HSH9W7y6v1rtfE07OyxUriyTEkMuzwEfMFQn6Ae9ZPRVsmtV0V
i4vRHPxR1GcNYiV8pL1jgmv922VirqZAGSfXcvbsf6MIjdZWa7dgKwUPgexmvhaMGDO9cVvF9Jdr
zTaauhYh2S/rg2BL23SzFgaSeITBCr3Ph+rurcZv+yQx79yqH1Bkf2CVD5bR+v+EEgOYCbBgeNlq
UTvZUQ5nqRinxpSHZfJzCM31bE9XWO31jMYgCF1KaBeain13dqZ2rx0sZHcD8ev1SKadfQhAEVm1
0UE6H4Neh4lMmmj9aB3VM1oMpalf/1kUy6I0uiMH2C47gQvoDj9kvwpgaTpjzCAfmuMGwPFNxJLr
TKHPNRbYUzMZjOwkIDTzabfLoU+epniJY8u6Gl3TT9n96qUBA6luIxNQ0cWg5poEhBOq9QQC4sLV
0PkohuiyGiqSS2HOo1to23AbKXrS9vwgEgiEaqA3WJ6Atp2EzUCGEBwopZJg7JPaPWFK+A+dvJ6Q
5s4FL/Kt5zpK+saWslHuFBtIaLIIysMOKV5azSdk09m56oPR1m3E2bBZNPHpt15sOtE4iK6Jpbsg
FD0FhOQMkbPDAnnmkIwvJwDTA+E+6MuD/pKG6YZ7hU30zBy63M3W2X7C329AOvNmbWMxj1HDWroV
ClEWq92RHwrQ3fipN8WEq1Im9xVzDg5nXU8CXnDbgzdkNiJy75XyGMoOsVaP2sr7QcxKYZI2p3ye
BJREwvRVl9A/jjKOlcnkOBlPI9hNq81VL5wSZvAiljST4zUr49Qon0t32nDTzWCBMhZ8lciGx/je
oUGvyYDOuXn7REJTDmIDkMuGOhe37PKR0izidktSVk2eZz3Qmw2X7PvnLmQocYZD28/Qcf9aD8Kf
1Qhtn6TIlQeTPP6UxW1wlt3kVWj0YuOc/WJwoJg3tPUYVrh3rMhPMwqCbWKvBjZTUskrvk0cbtqH
dDKtj4XHknDUzHT7Gp2uEgJPMn8Wu9FlEC6OWDIyhiHpw6V2mHILbk8G9zBMn4tk+M3hYkkkq1Qk
xEKq7+sK+3tVANvqJ9j36nEtbnTbLlBfTRUMX7Sw+5Yx4KCSUxhX4XRNpMKzKTr0hoMbnDUSGH8g
F2kxnz984JUEh0zAIIbotg9AGMEAt8+bAWHgdh2thtOHZRmvJBJZRqhlpDmOEyROnbcm1i1GBCRb
lQNbQMianKwTS4YOAsiR2vaxTyqDz0z8Xk7WbjQkZh4mhcWxssonPJkMtITmzxdJ2+E4I6xdFTWR
orn3cK414OvtOkxZuad0gcwORq4vip0tetWWAsrPLSe/KMZ687ZhemNgdWfnih6jNxByqh8/Xd0f
Qt4AO0VN4o025CuO/9DzinohMzzQ3VP82BuYKzynX283XB/Dplp/XRQBHchAM2OYelbaH5Xr2WhY
nAALfdsY65Pzb2RViQ7ZN6qWMjtF4HIB7eIQP+33TUveUV+UApJ4Z6RCY489Yek5v7qk6UcTSww1
deFx7XHxdBkdj0gZbmTitPScGBPM5GUQ/GYz+0MEROo3ZbUxcyL/fqzhNaSSo7hds620n2mZrOnB
xCsiM6dDL/r44e52ls95QpJiKwlFuc/vua1ukW8DVrwhP5w3T+5ardGzvK1eicjHidom9r6hvi1f
QQN1kG00V20g7gEz70TKh6sAHpd9icybyqsi8qwYtikOiH2kzMQel2zp8JzHwt4+Ka7X/qqM6tMA
IiJX2/QjsAPtg6mOkdQOEMpHi57aTOeIzqAMrod8TVX/38TA2KvwiCNhwsZSB6E1IQ4zDDNuHCKF
fLui264jIbRuEZYwFd5HHdZPAHWBzn5Za/3KkWoQ7p4uy0MHX8BVStskBN44/om9GuuBu4OSZbWB
7K1j7HJdvYH/xqtRxoe44v2T+IszRURZQqMeglbJ3HAi24RupBxK1smLJSeVoFHVsFzOfg4AMTvU
kyX9vQwiMJdBPGbDsBXhoZm/cSOsQJmNpqJpeAfZfklfuJOl9IBF9TKOC+ZhSy5Y0GC0u99rzvfP
otg8SMhkhILwoKI/bmHO8Haa9afVdrglyHvuRAW3OoULiITqT0nCQhxqktyPfzR/qkMJsRZm/WJi
s+t8PGHu/qds5c7EGlK36i7XD9pMT3JdPpURMe/n8Zi0na5HsIrgZBZbQswOK3JotSUF8Hmi2Aa+
v34Rt9ZDBFLgj8+Q33jjvcnp9CH8QMn/obA5Z2qTK89gfkhV8RduGH0allH0f2OeqCORB/n4RecO
sgr9PQd3UNkuEh1L77tXAgem8hDn/iRSM6Ua+UtWMHQSIiZA10Kjrz8aNpwVniDXzxyeZ/FQmTqt
ZYZuUa5XRYUJKKqrftQKfC6Ccb+/cNJPrc/aSCk4mDr1M2xsWQpqeZ9GQO0l7HGi9Pf7OXLKZQD5
lQtOInqGcHGR+YCo2nLxC8NySsnFySwOPiIyRqyTvP5KVs6r+RaJtjlo2x3lDZeswDmKhLDblR/y
qJfP5keVquO46Fq9YXZRNAgYd5y3N4yiv6BUAI7jeO4YOCg3RxofVaf59uwZYP5BCmDF2/pPnjGM
mwgpW7h7trlz5WbawtJcx88jPJxzytt6Kv9zB3G98LxG4hdmVMK1TeBnG0M/P1fu+apkNUSN2wbT
NaqwJDwIdu7hcpzBovTdbLwEaosNTRm4tm8EnWPhl42Toh9DUUCLMC5Jl7DTMjTCK2+JSV8Im69p
duSZaDLFDPud2CFC0JpwltdNepgccFot9NT7DJSrLT7IPU+2BMxXtWPuHNoqWwKztZyg91Qzg2sc
Juujy1d5aMlhgLBtDI3lZe42UOh7fzaqXA6VAxvJFqyHcO3B8sbpYR+6QWfelKHFPzyxP/kJ928g
AMll5DQAq9qu/Xji6meVmxBE9wqY6cKOPmM71vxeIJnxFUaI727C3wUza5F54X63CmubnMDQn8T0
9GOOWplguN6KuIQUDmUudgiOBDKjQLVavCC6ANdM9Z4PT5vGkMzya0BEhSP9iaPwcCMbt45hMA+H
xum2tru6CxxOafX48e5BTQG/r9jt2cbxUo5aCgpG4vKCzYFbh+5yYuu2bR9oBeYrp7y0qHIHgqKr
y1nYOs1q1YtQGfoGEVu95vaFObZw1TGM29v0LUcP37AVKMgJPsSsqo6DibD90owdKzopIg5T1TgP
+o3MBh5l7cHTaQ8j/ZWRfmQeEP8LMnRJF1E7//6ijOTnCXwsirDMTVKkTfR4CFMLS3CvgRxHSn8u
bO1XM4CTWYLh6dnYKw7ig7m03a5P7Ubmp+6D/ImDm4aLZ/IXhA1zggZKX20yfR3ARiRiiFHffW9C
iMrCB4jXd3YbSrgSFrvn5LddwS5g5AJKInxE/1PDUZUMWXBNVJ48x5XAWNlzysUnAHR3/EqxGriM
6HOvQnGAgAEZ1s4npSs6UcltYPQFB2tcrgim+nhqoTJ2kQISfbQeEcEojWg9L+49j2voeQxS1vvc
GM2icQuQw1nBhZbue6/WU6vpKkZyj///R/toZ67LC8n7lwO24zWxnz6lXEBbiq8aDAi7Pu6x1Vw+
SJTJr4FfsXOtx8RSyJVFQdYlZV42XOMCJ+O+XGsTkjou0U0qT7UyGGntwbUAEVqEpq4X/xhsVpXS
1BlEpgTWpIb+pI73QHNlpikgxNQYevx3Ts4EqtIZMB6E276GxvJlp3eSUzMWBBf0g14rBVxX9qWN
/w/c2yAqeJRLq3mF+MEZezAEbihGYjj+UjsXJ1AMUS8H6dwnPG0FLjccIf4r9bjbJpCCvoco3Ljb
/GxpMY3OVHNt5VzT3VD+Hu/oT80OMMcs5Zbm57cGoHq23Zz7Qe48L/B4ClafQu8GS6XbDCdMjzQF
L/djL/Ebc6tVtY7Jvv7chpjFX9TXKZCojIzkFOCw17gDLchX3ihX9e6m8+OdO01Z1xEHMPA9F+tJ
ctNjCjNzhKC5rUXrUAYx8aR//JbVKW+ROawyqTfskfwXVWVxp01ax/jM31VDFCu6WyhjK8LM9zYB
AJsiX1Ea0jKvWAvP3v/HGXit+flQtmDjb4FDXpNBOdYvvG630CcNcdbfZJr4D0aT2ltmiqobsqzZ
IT66sM/B7qOhoMkw0iKBe/4zVFsPwJNblM23Hh+aB8urAByE2eFs/ESzyQtvu9CNa+fT8i1p3nmn
MIqxfQiA1Bk64mAwLThC3ZD6x7TGAoqNywVzkIDGRrlNGjJL5pHZB5HM+UBgEZdn1Zk4yfMGBm9W
uGG+/sGAlr7GRhk4PeIa1Ao+/oz/8J4gD0N1qlc2SbfLTGTL6SRfp1EoQkxJuKC1wSUSoSeTquRq
xlOx22QnfVrlqSYd3kfG9Om7JMDpF9HJgLV2v17pcGM4BRnBd52uLQKTQVbuadGaSddFcUJ43lc+
0hd3H4j4ygfeJgyGQSOrGksvNiEINvpsjX7Ii1qfAX1HvxVMi37XX/LyKiQPUDbY6YGEfuexY0t9
cekRPEhf0daZhxozrzfpATD/UszPKT9A+kbBWHo/3qulk+SAwZVSwLq8/AokQDANpNdly9xUR55F
7Tes6LSe4Pq5LTFMUO5tyeIkoRTeobgn/Vd7QiYKDbyyOYL+BppOwdR7AsMf7GSFFZ+6h4QL5p6o
7/RRaBHf1ExtQNPetEBefnB07JHORUAokaxwJV6PYvJGp0VdWcuclxyt/MIWe6+31vSglHrw3cq2
R8vCeWg/S+Mbe00S7RvOl7LNF+JP6A7dk0MY24loH/Lv+2TmcQiKvo/AqXz5ediLfwSpK1K0VtuC
whgVITp5LlL2+Dac//090YyGaBOejycEv4B/a/RWH+9tNuYqTG8263x7+yIyL9I5RVcionpsoo98
OUlURPQmZo7Deck8DF1DAuenDkJvYHCQUTEuJCMH6cpm9M87Y1+RAQKbvDL1hkadlkf4+Xb4LlBA
uyjg1BlNs8GuTJguME/9IglO+7JjUx4dOO0QXIIm7p0HcDGsf8p0hkrKXBpOwg/ln1K0z4i7d+DI
givyp0FSg3VdeEBoFeHbJdu9vyUMUexMw3YfogvTr59P0sukrmcw4xuWkUexNgVNJVT8HwhyfjX9
Z9AT4Ccyyg6pm6x8ICTPI+oFapK3ox0TYWLAq+Hc9ftoVKcoxeQIe2J05b3I3w372GClxKGqPNqM
igMrHtSoyep8Em73f5fcWRq0gy0LKLOaXrq53ssMShap2poPEDaX10qjWO/a7TvcqiKw/4f3avkp
5Mga7Hdw98WrUfWtnCPmhoBxzhzE6D463r0bMOp7fS8Hsz9SXx92spzPGsD4ILSWqs0j+Db7BWe/
n7LZBJka5+hGnLu9KjQH/rJ0ubjKGTlaYlHGkn2jEYNyjeO7jaSMW0yTrKBQg5U9UEUrrhHFYzN0
DlIcZbg720xk2V8kG7hQNTuEGHSKMLcmPgEp9D43bvbt/viJ+qdHQkihIii0jTJcm1mq9Vbi4dwY
aVgNzld4I1aFpOeePc6HCDAp1oafJDkLrFk9KrQbA6TlqNVPvLu1xXtu0bvbHz7EaS1ahNv4qaej
t9wgUsmSxPozEQzPjFIR0DiPN0OlgblU7UFajSM57rF7uamzRKGY+XuQ7W5rNi4dlA7SfB7hG2o5
CaD8Xp7YyvcnHgWTIx2GDX0YOCydBLkyL6aj4GThrHPynlt52he+5qNpGRe+tvePFSNtXOMYJmw4
qNVV73bMRpCgABQBF00RdHmhwNtVf4c3kdB790WgfN9h6u2ZT66bQowsPmCFpozxxjmhXrCrx+eA
+5siBT3mGEa+xQU5Ty4wSNDPhBiEeQkLY8pN4tPT0Gxuepj69/eQfVd2FKhySbf0jqh2UlPhvWrV
aFKbKRratT+PT4NluXtpRRO6e08aCyNhh4KS4bKfWbRwgS3LAFwcfnS2YBUXScRY9F6lkwnCQqPb
V2JHAb2CZoq6yataO241gOiGfNWrDOupEB329/ti7QC+TVqIk6gJtrQNfRo91+7g+JhXlRRgJsHO
OKKk7RujkA9iY1RVvCS2qspIRiS0g/Oz7xNaj1q6igdNyu92AA+1kvnwUV2AqwQnBlBWBbg9UpPo
jUqa6yeV8wFKGbLl0NrzPK2hJS2C0saDJSp4pFUAR3KMH7PxuDnmjB5FLEpK1ikJmUHuZfbaOROM
wcWCe6rtQKRSE2M01DkA7ZxtB7VM7VP2Me9FFiQR1QoBIF3p5vccqElQP3mbMe0mm2ID7dFk1B0r
zpv1qAhbZCuQSDAQuicq1EefFWWuo3QjoNXRFfr5uecF5HluMlwsltr9hhGANLKfGSwFTxrmRsYU
xzEbcRQRDH1O3svNHHVSzb4mQ03QmjwT+ppfVns8ujQsTIBn2CZSWCForYytICSKmBm099OOfHv4
OuGtJl9xZ1Htp39yIWHRPmehB5zcHJFcmtgO0UnQxkqLgy/zWjfYe7vAMdpWiyGQlmkFlq7/Wagl
6+LUiguMiy4HV1lUZQzqnwbsXdoXdDWAtHCyGrH6tj69FThvhUixjMFVOsprlkdoYiguZmTbbo0X
MLW46Lh9ce9NBWJFy7PXimAmjM4i56xErE/5zVsyf5Qh4hjB4vfjSmf55R3xdUP2xZv4ZvO+9Olc
zj2gW1knlGVo6B+JKa6JFUfrBgPV6blr4BiifdYv+fBjCdXXWPIKNk/aVzd9zhGQHk8y78tHD1S0
7LcjRnSgiMxahsSO0PDtSxAOm8agoGwI6h6B5uKyiLy3Us1CSKtO67fQ4QzKHqn4u7gApgRXBdfE
bvqBH/qpy3BqKHUxknzc6ejpds5ZERYZ1SEROkdkTDp4upGLgz+gGJUIsjpNk272NU3suvsPkpj/
z0t+GoIkUYe3+rzST7poJXzAWQ0GkgXa+BqulCL9Wff2DoHHWX54heSFHpnl7MnHwWdmEe6zJF3c
b7pgFOuHurFN/GQHjNolpK10Ay6Zor+u/12ExauVVOms/RwOqhtLZsnPSf5/BHUMpHM4WG7OnSeu
bZqBPCpsCkcn/nxadgbOHueLkIR6Hper/OBvGXvdVoSLbXit5ntiyWmPKPuxq1EAnT7FaEolEVII
xrUzOulGb2F2lYnT7KHCByDcTz4k+SQovW4Tqc72pmtOupnNBdKQfzF+b3g9rYUbWTk2vNlEhJVB
9yTqLVClgTVXgQZ4U1CRg/m0VSu6/853PTbJb8ePADqqxjEPm0uUf+EiICN5rUgwKROVckr/FY8/
TLf1srqZg5G93bNvIRflLGCVlspugFAo8M695Gg+ckGWqHfM5qhmsM5tgBE562BuzaNOTZKM5oI4
CPdp2+do9vsIYFY19+MrIrptx+dDHnriKNaa3Piuj2q1uDBc92HSyOrneklo3+Jtwz3+KPbdYdm/
vCnYeEjPZzI4FjAMuQrva3FWxmynzkZomh7WTlvGYMcJD0sDpQgwqlVyKB4ysiehOiNophdHnMAg
MaeLRPPq5zl51sWKjQv4LVhs4SHQPFT+4nDhK3KpMWD7UaWAFUjeBU+KB4deWwj1qWkO2CrgleKV
ja8mBzaB8Y8FKohfGRDBIEqg9U+/aiTqc1xF3WSlLfj4lLHbdOahp1jrxmTN93+L/9mIpQQsX4rS
rjaxPI/CsKHmY0St+Ie2kgcfIxgA39b01qVXW+VrB1O8CYxEvZI1OwG5kInxx1cDzXtieOAvXUM8
/QUKAF7lycZ27hrRlSN3zTJRD3EJ2ED+a+Cmohqu5a4Ra9+sHOA67RQWUomppBSeC/hGAb00XglH
T0/8MsUFz9znD6e2KCyO0+COVeA5IOLhW+UVC9DRccj+aa9v3r4JXW/vnIaMqO5TtMWW4FEl26Jw
o4x/Zol+Ueo2Ie9R9TaxRGgr2hAaH3Yh+DhQkaScvu+7tPIhdYwYXugobGSTcUGJm7xqtKLm54cW
XhDPVOiCfaQK9Q7Rz+j7VLc4VtYwHhsJzAj5CrEtbXz9vmUYMaiG8dntPO/V0fEdUK2BAzNbL5i1
nEIbMUyMcwFyXmHIOvGFTSpX/qmbA/m78qPj4v7dgUsYnGw5I34IBerlWn/zlDvjoioe2pHsBVKI
zRtjRmuJJXDqHbSXpuWfHmiJ4U7jqqGNjeC2iTQLkTlet7hhC5FfxA3iPNIIoDTDjrRrmzqZhPvA
ugIHwHQn7Vbhn2WOJsNZsZ/30qebJDIKuyyDMnhz+1flXylr/n49TaBxLvMRrw2TbaK3nlRacuGD
rAhBLbuJblxTtamSFdL2XDGsF6LEqxRIxblmWEcQznlrSEIAmzfKka3jyPhkWHF8fCYOqnPNMMXo
xnPX3Wf+GISKMBKlynn3JkngRoyvDvONEPhV/UaV/PnxU9P4fSOFNHQnXM86wfo/JjKSq5Aalfh7
/M35lC+ftMhyoVlfgYJdVRE+DCzabSrsiYGuG9z+bC8uUvyyIdFCC5cqrjmRGq+eTddvO3PNn8Ql
e9q8Dsy10nNRP5S7i0Hlw9egb8IrwxSP3L9AS1idIoowZTCzwkO//3NYv6qiQY5H48WaRmIOAqKd
LB4agq0nXY9/H7d8sllXZpk3Y2aI6oMAGSskI2stgNxRB2kt9TYwWFb5/mSArNNoI0//2z4/l99/
4Cgm5JFW+alaMtgnbXgsN9sk4dbOb1Ehgne0v/iI98P5AI3L14/auCThQXVPj8kg0PPWoNmPBgMF
XzT513WiO8NAbCEOH3RVGNxT8MYahWSQ73lSAaioJ1R6KdUbRczcy1x8vHqrT5v2ETMaKbInqIC5
xVv4xcJxp2XI2uXlmxhOo9jlV4UdrnohoTBB05L4xjZKp6TWQX4Nn1fwLEqzuyrHE1xPYT7twUEI
98ahNEsKKX9mbuZtagm0Vy0gHR+ra3PUGnFbe0nxiLDLd+wSUWYv/kBNM7yCo8qjOsb7NyaQEORt
+udafeNLwGUPPqmc+DOn5guT/WlSFlbn8sCcIu1R4InLh2M2V847riKTsHq4qCO5l/PvZtOJB0ki
eULBbgNO+0wN51Q/1y6EyzAhgDOZRR/dkS0IjL2jLUgRse7+ABiROFBlNnttbjiQiGnEsp0ITfw9
mFqR5BRhMSrEOqO8KGYpsDt+IBH8wfhUU29I29Iyab+hFs9CYiP3Q0QQmyBidHBSoFxXZfH4Xg9n
SFWcAECH1QGSB5532ulWKUB4H1VnvcT/FNfP2ahAXCLa/s42NG1esqhQfQnUR1ohHHYenzw5Bfgp
ZSGSbrmYcgNaPC0zImJW7Vxix4nC+rPS3eTz/27SRZ5/XP9a1G1gRPGfOyLqhKCu2l60hisLpLU2
d625j6kTDi1FgWF/DeJqC7h1sViaBi2IFRPu1bTO0cJj7eRx9h5YOvCRGTxPS1Hu2tLoVBkkoYJO
x8j0KEctrZXqUfQ59i4Pnjb2wGGxF6RIDWrE1N6px1MiTahmPPryqzlHsms8x7dFusIz+mX05Bps
PM95bUlRkCJuPVmxyoK0rIuwF2gr+Ur2UxZL2cj5vLZNocgmxhjbLstvoGj7ZVeK2eeW8Qj+eeLo
hxdW43pDp+DLLXSqkMTNuEZ8459zh10bs56xl4ktNFMrWyVDpORRekLg9Qd2f4yfNyiY5e0dk7QE
pAcCYCPTxdjrQaU+0Xdfukm0948AXK2yOwX1cMWlWm5MIXhR6RYPurCUBgODSeoimA426QOWQdMe
RB2HIw5U8UpYXk39r6FP7acwTufHq4pWZpa96ax0skZ6wD+eJM3Iw+dG5UdyntpDC2hIqmjXt1MD
4GgkBCLIV2hO6CKkEFIrva3qU8QxPgIQou6WAW4EClXiBFNpLGUcJW2/MLcAOlFiC5l3TILZZt6S
pjW1Y50vp1XvobnIKHNA75+81Av9ltNoHa0VPnbEp8D+F99tw1NUj3UEnO7zz5IQfJ4CktB9UV9l
3QhVcAa5GzJurJWEfi5BxNj0ORe1VeapGLxWJ58I498Ew3BeT/o5b6DK3xeTRHZfoc4ypzysApcZ
JqbcaT5cWg/nJGMSsDkX1/6wFZJgxc3xyneb+htPS5YAke4DWSmSlBeXekSoA6+3obTWKUG0LBab
xHdoSTckDAhNxi6oU4g50ga2oX0yN0VC230VNkEb1JSDBBucCTWdzQk+ZkzGY/BSKMbEK3ivDoa0
ZLTE2vEDf2Njm47aYmzCx4y53/KJeUfSYG+j0gGwpR8ZRFU+LRFCMId8lfpOPBUiRMfa0Ji5LBhk
VYSvw2+n+VG3uwnvz6JBBg4lmn/wz28D+PQ4XVRMiUQqZrhFdViJPtmWq8g4lP+yTgnbY/SmSVWn
tvLC41xHLq9XsCPrMf3HbmL8ua6OIbCCxaAsZCIoSjG7ipPh3lx730ZzXQ2qKUdk5XyaVBLuyM2Q
lJoUyxS0mdKIfRPuNNRKB1bqPDSI9l5t1QTf0eRtQPoAGdi6kuugHfe5cHCXYJdcmATrnUsDInwk
kxqh/02pKZ1bRUzGK/8O1ge6LnSBdA+13UN4AHiHvEgCqXg5N9aaarpPyWZz8BtXAHRB1EvbwI2U
RF14qRR0WmjJsA6BtzTThR4ZAsLIWi9Y0mCvJUhR1EbC1dqCVUxBxKFJPauyMljSNDyssd++uiE1
bNb7qLO2uoXqiOmkY2vkN0Pvliggdv7MYusCP2Yf20bjARN2Tkojxx+udGEx7K35F2JfSqxps3za
Zuvy3GgHSTz305PeFkGUPNkxLTAs0NvdXryFLdEjAwVVEnCZjUOgSSqKUc+8IN8CuS8ADaJnFH3l
YE0r+e0B/FFmbvxyP07SN+bi1X7FaI6GP/Q6X6qXErAOzuwRuGiV78NKNZzpE2gkMXTFjjQgBN40
7tbb5d32YtrI04nuuzR8hetsWFHX75iXk9F+8/upVy/G1M+kwgs5tnF4mJd1Z2wo1+b4oEp5T4Si
pBzHSVqRH475gIvhf6xu+Tp2sDb3f3uR7/pUrMDaa8ViLLS+0xi8xcYndrDI9Lmoiey6434jEke2
D369+zJ/PdI77v6ESyd5qQEM+mYI+/tUsrLm02xoEyqdeGhaeEgfdzFrFiTaPKhJox5d471A2AMv
4EvWBvC/HeCy8LXqmDPV67NHSg/d/1CFQajziu/DWHOAK1a2xRrZjk+tuGcxdgd7VY7eCm5H1WY3
/6N4kapShWjdtyxAXNze2kxFL3s+okJBPzKZWPISxJVv7pJukBNXdRJ/0hHR2i1FECVmaNFK+KIt
VKsYpe42wFHCB+GgSROWLi3Fb2/EBeXxjIloPJ242AeX2VYCtZx4bCAYAZZp94Ukstqo7NWDTDOe
dj+LvtQsED8Hh4mZLO1tvUkIVqOG1HKfuhrxNPTWzrhQLlHNjaSkubLEQAq2Sz0yBp6vXGkeUB5k
eEaG8KFkCwBFJ9hUGriVP8CBY0YQniR3NmSVwvhE2vpKaocFb6URmdkrHMQyszyPyKDuNF52qMDX
oP6LgV4nlENTZTLgk5/pTZtFaP9A7zgZOpj0lC4aMJiJXqc6TzMlm4XkOmflaZrA/1j4PKlNAy83
nsqy/Hb025QEQkpMLMzkAZDVuYe0qdOj5yb2bsl9nTG1su5U+LkfRa8FL3wmDxvDv4izBmydMShw
sEYywAFHFKNziOt7ozzCtEtBI5hu3UD1Ss2o7ofdD9k4s7LiznpI6JaBpHSsuaQPdK7VgCRLmcMH
LxwLAbmSaqhpg4wDicehGxGppblyYlLhR2N4rc7N2o8YQSXSXUErnvC5MjjRp5Pm/MnL8hjFBLy3
t62NW6p5IcGWuy5LMZ/ATRGZtLoJf/b1OXq5H7pIHfgLzjlo3WKxT22y3OhkCOLWL5Hf3Dy8N3R+
uOjYwdC2gXOTjyCqWRiEzIctGEDFXXgvKIrQ0qjk6klr2wUE+cV7r44qk5lpMNEVErJ9IufZaa2I
+/oQosaRJnXyD5z6toj3T5g97mLT3ed7J1kxIF5cihKkcFcR+6Lydu4ojQr3dXB298BJn3SndYIx
VMxAfOUb4Zio+DvV/lH065El9Sd/SrePXJ+8ulhm/RLCte+up/EGRxfWsQRFFI21n6SwFx/JlXE1
HwV/rAfjxosXoAm+RpkP6/lj0uwKAWFi5h9QPz/z4ZwMWEtir0jP2eBFB5bmll7UMMXM3rn6xv5w
xUuiqVvGs0sOISyWI/ZN3aJ3euMyvzhCDYy5X22k6CTBVGmmVnXDXhJ6W07P1uw+Yei59BO3rKpl
ZKyw4PewxLRsmfkzif1DGvRRJUMqx8yKgkYD1sGgYKThxy3XINNlj39Kw+H6+ovABCtkFl35yXbz
gAMU6VeZhkl3MAumm/46yqyvEsAtL6Ua877OfR2/W9+KfnU5VrqJn3bT0nKbKYykz1FbRNRQgGrs
7c94dQ20t4XkIRpGiRr7GO5fneqY9p7RrkNqUQmdVyij5BKVrtCyMP0ME3ivYJGqwmRRBdjm7+vX
FggOUDeouUH+sBjVKd3GoAwaVNAjan1LpUAn0f5yyhvanF751lew42vN4WxuE0HDwOADEwLWER2h
89kM2pvAdkeO1se/wIcm1G0HOvvv7AgDwhqCvMfW/Y60sMxMaIbRwTwIbryzA5mc1QKTjEl4m1n0
BGUx4PO10yEjhPC9ljVYTp4gekUyWm2iORFQG7RBiZqLqdgUeCD8EEm0FElt61MmghfXD4JRkhNm
jFgT+M5Kwr2xSPCLYaRfcvKB+nklEooBFn4rJ7oH2Y/9/mtqbrT6oaMVb0Y2B4xOX+dGN6JnWgNH
yfCqwur5p3vM4qkC1VfUL2u52CkRQUlBvR4yiPMy7FcfEVjcdmsV+IyzQF6inKLjBiBqW6x7gtiS
CbgCpm+MbYpK8nx4QQokeE1yjhYxSfvUDXS+xnxWEdwuaZG18VeVwugnLdIhBzvgcrF6nPQXyBu4
mqOn1S9h2ykK6HQ+PtQJjJ+eFFoXzcKMjWC2jGEAVcg7oqx0gAKH0fsAkBn7dtej0p0EDVJNY5IJ
w+Hi/LNoLW6yXGw7NIhOkCdQDxNO2KZTcyiN9aBz3HnyDZfSo+Fons3ocT58amPfxTntRLkZHg9g
2VmACqqs7M/WJPsZkoLcsefYiFNbw4LtgJQ2y+Hfbgjmpsyh2UILvfkzra3o7/7V8hc7j6rv70wH
ObvjkYGuerWJbrnZ13zRtxgTsXTd/NKIcGa8Gmbow0T7wvA1MeZs1IQKcSvjCXtd/VoPV89ArejE
Srjt3/+1+VH03SJV6RrnV6bcyaLHVtoKUl9C/TmecO8Rk7ravPvwaZkxYzYUQjDG4aCv8gPZ4Gd4
Ij3zUZVydXyFlmAuaEoO7xjz12n9s1O4DZo68RwozXHb606OV41dB+ACWidYuRqTdU1P7AYiohNY
zOmtydiKKheHXjLqB8xiWXt21e9bMs/TFqQ48EfVuo/33BN2QDR3WH47cWWt8fdXx/dN9ZgyjFmU
1WoLOlMckunEspoRajrnpza1aWOqk2k5Mo+6Qvb57fqtRO/KZ5fEmuZEkdEo1R/W28xxcNPt4xA9
QjQrsYPXoF1bHRrNWNI4F9cl2os7yhRqaaLkXCgLBT3EuWAfJdwz2kYK3/lMkVRtYD+Zc/G1v5eT
0/LwJI6C8quzZJAhznF5mIhB5PYfTBzGCZZVAId5v8Z0baimy91YL97b3KP4VcXzXduyRcWK1r9G
tQuhIANIP8CEzZXtL+UHQAPFingrIbk7rNT398U603xq2cwsvhrZxqNAQt7qIVw7huCthrw2q7oe
pYJbmmyas/E/44hUP3bHWWs3mlBduDZBoZBvlpCIdZj3ZrIPlHifHDQs/JE9YU9DkUZ38oXICBeL
xHL6pgIXAV4tXWqfQYn24QzC4nx3a/EgmI2sAt2gxOb8g7PEeBXMEyVPCA1+TOpfRFb0NjpFsr60
HDUY2LsEGOwB19gFIEkSodkc2e5YAC3S+I2qxGknXDUCCOHhtOSZF1Mqb3WR5FUBxhmmfdsoEoUp
uBg3Bn9w37X7uQQHVJx7JqZ1qJdMX33ec9ZQvkiUTqeBVW9TbvYTL+K2wOUSYq+nKs1695PL1G3s
7/1oc0wv/A2vIJF86Juv6TRk7FzzOgEUgl1vUzAa3NFXCKQSZ9P2MC/hwz8VE7wVycFJHyjmIDJl
6M25n1yge0x6DdRrv1FjrMlG4TlCEabWpLBqerZr3Dqic9eI1Cjft08cd3w0cVuCnO0J4cF2OMVc
uv7V1JxQyINDUtlvrHsUR/xzPAmNqR2UVJYq2p96pCT0agbq8lUFRaxaNplZ2umfPkopvQPhY8jQ
gMbI6a2J8+N0OzIVl6k8AJgv9mr1XgX88A0HZ6FGAcNLg/RBLWvwNwrrrdIomA0ZPVeasOzM7mKI
Ag5pPfK2Og21BOSBTZ6BTxuZKquhfXhgqbeoAonThQ2CmSPllJdfP3cHdYQEzPzZPV2H3Q0PBavT
rKOygSA6U4JTv+GHS+Q0qfGsy8bGszGaHaY/RsjuUOhlR+yJpFHsDT4ub5Ci5G2A8i9mCGgexQog
ewZdflyuplPdWClgxLvxK5Cxj2tmpOxGMjmFmavP/RLFkp4N1S7dspyz0qgiCEssRGgcLQDkNBhi
d6/ht2WHTMkvxubxXn/00lSeS+kKFIZguY8bZv9t29jwdQUOy+g93CrZ919fAXjPYr47DssjgF4i
l1Kqye5ia7Pw723YQF1KiG4NIyxoSppGBmczvPU8VQBFww+KlaRTk9J5EImOCGvaKCRCMbuHd0l6
12xD5qqeA3bOKhWxiXBDsc/hdAOyz/c4/IfNfonXgwS0wMEHBLVbNjtl5QC+olVeEjV1VqqnYpcn
n2ZGA0oo3Cwia718hCTzV3aVcleMsTou5XP9l0ivAMW4rhtOmGLABeD1REVSI5cP5nuRMHsGisjK
Ep8LK+O3L08a0hOTg4SDqns7Ke+EPz+oc1Ekrp5BBvqKBEj/T/EAeGzOixfEuGsIpR2+opZW5+Q1
jTu4jAXQ29qa6fsF8kfp2Z1T8bz59C5KpBfVx8vwugUmv9FBWHKg54F0kmU4hnE4Y2m2POfzsf6E
6tOHlC42aWkrOLrD0g0oCanghTkU2A/zCC0nRFyw1P+jmKQByDRptelfrv4ALBOKP/LY9P5MiTAR
Ve0Wy/SyyccoNLCTGdVzMEagHafLvQn0nRqBU8faY/Z9GDAJUmjDbyIaa6ec/otA7ISZEmzr0rlu
TXjpNYubI3GH4YBPIIqdWrIEbvlwKwYsRTEjIUWz/icQmbZxXJRlHih1KqegZncMrPK6tBguL5AZ
GZa63qI0avIMi9lWj2KY0zz+d0IbgBGhNXxG8rNWkb7kewHHGE5Pqz8qLtIprV15WNQQjCVxC2Vm
p0IQMt7rTxnZauRHZxNhKE1XzuQ/NtCzkCqUe25ZfOcIYhAP/f9cqc5WM5Y7ix4YK/OM7NlLFiyI
WhHuWSksm7hkNgNoj6bbQS9doDwsM5YKoMRBT9Uk6iq3xRTGNfzmYLAgGnjDhtRD23sRgOQMIx+1
QguzfBShtHTuqJtaNEuMNmJ9JyK5R218wknv4SOlerYSJdBa2VFPw+4hue80zGCjagTCcH10ZzwM
Qof4lzQ8Fc/sjUxefjPcBdsBbTrCkKdqCBDNoV9ZmuyjU8wSV/RQxanQr+NJIqSxyF/vUOqWW34P
ypifvcS/Xcby7eokJ61r8KuPmFvxY+1a9NTU9xL0nHvPag0pQN8enpeWkxwVwOpN8aSWdqFznAvE
yfw0o499D2z4Dne3/bNJ7zMqIohFgx2q3c/WsPGtTG9iWnvO9OxWCTJpqhQ2HfVg4RunVLqdSPtl
7nuUs1ZxkJGtT5VC3i36a+GoSN/wVu0jULSuMaeMSdzc2UJjnq2b3pad+L7DYU9RK2KlWMe+l2Uo
Pssem59oieQLs5jRztAkwqJYN3MwK9mHKp/aq8ErFb/6RVKTXOPZHmzK4HGPSGV3ULri3k5KVMU5
53aXX6EqaWxj8Nmt15Fjdk9YLJp2rlm8kHoPU7AESOE5nHi44yHZuv+IXD8yMvzpoQvPrFQg4Y1M
k+fG6/r1KHMiDwW0iwJY80hwqA6nstEs0EamRFOfjGefHb351IW1/rBsAtZbYGmkIOgT4zvUuA4/
lFUA7DkniZcRKi3YsF/2PGwXRLWb4T0tPBHQGkMIXyOPGAmz3IiiJpz13xrZ/fV6S5joo/zc0X2k
hl51dZuH/JEHJUB4BelTfhQJBWPfXH96coTcTV4KR/rB4+FTxw7asKwfktdtd4y8lim4WgFJCOkc
/QUTCcS59kB0GAUx0Q/3Zp2Qrtl9XGiuWtG5ALwEOlueST+RslYE/m8GpxdRsoTYft7us55eFgzG
4rbdQogE4MsB2QtobHAzUYn/cJ01rfbP+8lQ7WiftA+oxsT/XUe0P/LKcrOC7M1fdoZ2I7pNNQhw
qE3T38Y2ndGWX1J3ZiJ5PO1WycofqdkpOnz9lvMvKHPdKww3EgW4F4GCvs8O2/i0d/4IKbKLxSdW
mN1I1yU8MPJbUlJl3J3/e0nn8SOV3gddMvGbq/nhn2q4EHbfcsWE6JNxmhRHi6hnCbfv7G4em7qE
mH5dNOPIkDcdJ9vnzK5gBvPyPkGzckWbQkKxULUJDs5JcfnikayAzr+1U/ousNOSKxp4Q19+w7/O
XGada3/BGOdF7rdlph5j0LqZFLBRp6MKpXjykhYWAt8X/Si/g73uaZmijOAB86eXIW9MkTogfrry
k16TxwOT8VH7JV86POSuRjeS/MY0Avg2/QziF3AQ36zZry88sIRd1iTdRxLtG0vvm5PE3bddSktl
kkuKG9Ps5ktZPegAmDdSJnFr2MkqjfVNBgU6HmyFiF5jhC/oIy0vyjtTVCFcKdf80uTZ104X+gKT
szmubYSU7ROREOgr5QnfKepidq40Nqc34DSIIlAx7oLXg62N4TIf7XjyJkKBm4+b/sHoHVQvaGJV
Qs4xa9P5coa3heHPo12J0l7+2WH1oRVw7ZdUi32HU9ElExgzg+GafuRztdo8WjungAzHjDJPSWGA
HIZp35FD3q1sUZGf3WTwcJEGY1CKSnItz/3UobTxjgmR0Hsgp3+DxbRLYEA7cNnavHUwGRXG90vj
1MuGcseS4A0Gfs2HpkVecuT/ocLzMTs2+QMTU3mgLg8PLBQRkz2kiIf8GkDAZagJGi2C7esSk8/u
zHzsaldtY3k+1Q+T1MmnDxI8D/Ktlkm0SwPlGEZpxOWOcMQZZzN0pNq9kb/eZV7REGcr7P9iOwQ7
nLNb6AznSRx1rKYFq6OrdeWaJ71W1D2WfXS4DWl8rO9gCC+pGKIVp0uIWfCL2pNARvV48ChjXyBQ
Vu1224INSSTcWp0kmSWAKMC1ec4LEaKh4Gjb/I9JpUZc24raa4J/V36d442sr9xDfiruUitt4sXu
Vd33dk9V5Z8AvqQ0k51SNpKSrfW35nKtKIo7K23/ql/DKpZJNiYpfAXRoIt77/dB0LBxdRz2TiDt
zPZuR6lQW4cVL1Bu2mwU0tr3atW/VgfDoPoLajnqFp5PJMeu5rxaLG+Md8gCQ1G0zuy5Hl1xC59z
Wa0UXyiOGzrfE6rpJCm/bv+3y1xpqa481pTDwOdG3Rrf50pLb4IkNfvXI/Nt17CB4e+oowXHnAm/
8me9aC29sJ41+83gXjUT2hBDY1za74fSsXwGSu7hXZMv+r2v2zxVAJ3pVMNHPCtHTrqNL43rxuYb
DSn4byBvyK8WJMw0sfbIgWlbVvE7x6wX5yf4z1WiGyLyD6dR2C/AGba0O3aTZmqakC8MOvStB2kO
JhOOeSIH6IyQGaeIHTGdBHyyOwQkN8Ih68MAz1qP2XflynZGkCn2hG8Of36Wz2a87Lt2Xp7OUOK0
YpLt2bZ1trGyMD3gpjOOWeVNTxpqZ3HBE6h0D3E35d9N0QS0TCvNw00beia0Te3JUH2zKGz92HPY
LwmP97LLnQFYMtxmFlgkvGsqajkCzzG9SKIAxNnKGZZH8AUBHG51ARova0FmWE0zSAL9Zo6TAjFn
CSpH+rUhkWR6piyU9C9rHXJC9pAvZvlYnrD6JIhta0f2TJzdX7XJ8RhxMIWrQmFAIfEXBn97LLfM
1wRtOb354uTOxySL2UE1PjBJevQ06TTAAH9W0b/tyiWqOOEyoYru0eVkgWrPvK3Q+2PHCIHaMJ9z
jkTQFkoMabnTwkHLRmsNhVO+GZ1N92iGcwfKWk1mRpZgv17g4TtxU5g9H4qgKXrxaV7Fp86kBya+
K4JApLsaMp+lhrQcqSud+HfjaXLxrm0IYDZyTUH5Ky1nYIuzpHsiM7dsnopOgTXIugtGN185Fa0F
Wt6jlW9UbvkRQtlkzv46HTvJcb5eUVjxpjt2BgquEYypXfgNAnIqSJrpVROxWShC4p0ky+dFp9z0
so9SuQFKw+25/yhFCAdES1MJP44VHfwGjQaAYvB6umBppLfzjGn52EEOtVTzGoo7vyjlpXdA7gti
8fR4+919FhwedcQhx1f02dWrXhKSyLw4/FP8GZYCNno8cSucOGVsxJNodx13WcL3iwd7rt8O43rG
6z/d6+q/vDryT9Dd0Ij0ZPpzISmxcyurPzM/HStomLnTDmBL94IQiINOxQ4//P4hWY8M1TetW5V6
e1ppwTWHX+QCr17wVH9Mx9G7zx6EuTECkZcLmxQyFiI6P+4JVTEUnczjyzM7nQFbpWnXH46O+Fuf
CZy69xyS2rUZ0BhnH6twXqdo/QKsYPRT+l5grG1aCGttnHLLRqhH2VsD2apeUiENHnRrakYrOB9z
efb+LrTDz/SrpNJlIrkgm0QrNbK/XIGjU5Hc69U2c3ytGvsFCFfy57DwuAdNDuDuv2cItWMg3GU/
k28giKe+Zo7n/AqSqf8Wc9aCo2WIgaXVwrr0mmAUl5hOHiCZ90hLv5E/0SAv9dYiqbsfHrq1ZaNM
ZYOYRqzigy4HbwkHPQkhKms4C+670xzA6YHvQ/r5EL77/qk5Tl/L8eRKViKLGVZo35XXPoq19aC/
W5fWoD9Uy/YurRXGIHou38D384GZY1PTmQ4hQGtwAhPXmduBZAmJ1Kzzgrj/8SBM/1qz7JJGZLeW
m1Ned0IOKF2VXVNW0Z3mypcAGM8ksaRxYfL/ug8PwQZnJrANtN8nAcvNPkwUb5IK/0h7DInYBBbv
TEEFcsm/xWrsJjm0u9efvk4cqzrfkVtnZYUsMX2Z5FsSAZPuYtEpNYESDahrGQusx5eV20/btkZZ
FEdZ9jie+6mHlW1UDjD4I0hrcGGER9NBOfX3qZZJAj8VdBKeFGObl2HM7+rYeQclWkWuEFBYIUCR
MjCrfLA68tmJ6hqAiE/16kBTuFXDmG19Xjlv/kRGu9vI4rli30lQ7KmJCR+dVYMAoXKBE2E4ayfr
rVTBEhoaPTS9VF1mYUk12Dhd6xlNOEilyXzgkuJkr/z4R0RtXTrok9LbAqqPqIWqXebBMkX9fHAZ
xtwdymNl+lUcGVtX+892koCWIW7rv5UDqTAYIzmLwfkzgkLD15KAVt4aYLthxirbAY6tlN3C6n9n
jHGaxorxOoIiTmy2iaq+93HH5x7ReJhc6RM+u6qpvj1FH1dw4LWeNkf0VA64DTXZiGeF/BxUMwrr
irnFQIuraYk5glpSJ28gvCFK7wLg9y7/HNTMxW5pG6L9hEWkttFxvkfBgjqdglVpA+OsV8KcvPr5
R02wrHE7lTxIH7HFBWa/azYadn94nnEJS5dJPycPxbaRslreQoQspm+483ZLJi/6CaGuEFKdabY3
nk81H7xf5vYCZjJBJlSaBtnjOzDgZnUJiTNYBTFi7hlPrv2ZZe+ZOXAbJoqzWT14LGNuuunlVCAU
GxEYjg77fy2+w4LtILNL/smFCCwIAF/vw4Jbw1P8JUg26A42MgI04DCKcy2Vm4t41GbdeGjif3Jw
U2cVnxkBM43op+1FvXIH/cgua4oQkUieQIIxjlPm73yBx3WmxDQ4JZSmzHY2j6oWUIFD9jnh4vl8
j9YQKf+7PskowhM0rDJERAHjQQHL2+WkqOQ6sdaP+aNNtWP817ybx2/7078CL3qMJJ7jwhwWl5N9
YzsFYk94hNlMAS0wBehtY1RUzr9GVhiLPKhHLYJ3bt8pIdFaAGladvmUx0t2x8CSQcEW49x3EoTx
My1417kLHnVgumS/RCcSA6GL5s1L2HoqzCY7NNgXGPlJ2mfi/kruMDZoOakPoNMA29YzDJikZVY/
cNs0ITfZwCI+HkPMq9MftMtlt1FsgBk44eKM6Y16tF6dc6Q7g5YIZAIu4v9wKZZF1kWWJ10jPyvM
XuQMOi66N6SVkR2kBwLDSMx6z3Dr7UhzGLuIJ6v1r3GXqbGg9iVdVRvED4X1XEWERUhoTjmmDMRZ
qKYtdbfREVGMG9xDBW69PTEJEDzv2VNgdaZj3BPPr5wFCaOVx0JZtAgspjqZ+HDIxuG2tqlSXYAR
g+YQM1oa7u485LBqOwWG3ImkScVnhOSBdcufNAUhSs7wfc7jkNmEJW1eB9AplsXPsGNCchfAeAq7
OcPK+EzYAklZ13Yt4pT6WuIBNwqy0YA0IU9BDwp2r/y3o393D13PN/i2WLwROuxqDffug3yJFI90
/uvLjbOSZHT1T1bYtCQ8yfrEhzaLgW+ANX6+5ELdAlmDwkVVQE0SdhXX6S5valFG4AyIt0kL6NrN
51Q32/n042sEdhp3Dp+37qMUFPvE1VIlQsRcXtMNeUwAPHsJm1KX+Zn7MYz/Q06n7YO/xCqc8gMg
ldfFTe/01wiveAM0ATxJPOKBZSY8ZmaVYBKM4c+Bo/xaEGheDoh+528+NAxClXaWYC7HyDkMHeAs
Qdtqgj2xC8w/g9DovZZ3bRyfFzmMY78F27bBMT/LVuZb+1n67nFEiehg5HDF2lQKh1xbKAgLOTr6
bDNvP9lTEibRyDUdk5MGzn78LJPsimMDcBfop0xFHvXcGkepwOBa531eTWA5pCGmodnwBzVO2c19
nWtGhPS4qlfXZ4QYyAKJnrRpRJsQgLN9cvvRFhGtrQEupnY42US8VoAysok0m7Usg1O5nG7uWQF9
Y/6I5nqg/E4PiHrKpYYe3+W1zcOrg3DJPEJqHZBRkTslypkmm/MmMocoG/nJiKTo3spCMj/RD+4Q
sRvHdBRMtwbIxjX7rTam9ngj6/lA8cKwcFAvtfmEqDqxpo69kSsI4H/s2a64JqthL+BWIOvMvWho
ueIsBRti9/B3JkcTuG441mpJlncyZFO+zpxUXJqqT49O5SWBMyHgJMy3oqxS1kRGl3f59WEzxGu3
+kS2zMToATVm6FpZ5b7M3vQGoIGwOBcX+dPKdc9YreFPmMKsVLn+TychSKuFZFIVLFNWKBGRctd/
R0TvHWztNd4Iw7YSAuOmsBdAsquNkZGt36CPe8xmwXx7AiHBNGR7ahJ+TPBSx9UjT9qjvwTvbVYR
YsF6m5sTYO3Ec8SXmXiREab+opNRVgd1U9wxi5SAwfNG070F916Q7miRfb0rW/k5lxcIFBmfZRQK
2VqtOoxN4y34eItMUsRIukw/XokmPoNhCO5p/yvewqdn3poPamROMxy4iMfjvdwAgPkNVjhR/f1T
0HBAq+i4JC6BfZh6+e+AbJCWjMSJ95vT8q0jGY0wN8tWA6SL0LVUlBs7KOL8fb7UpABTbYl1aGTN
2EFlGnRHhzPN3l+qV+gExqHia7QqKZMNfWa6m9fTZGumjpvpKURY6habZ5RP4wjslbVq/SUD1kVH
gQLAK66zo3MELEdZOgbAG9MXpYkQI6zBT8DY8iKZzEbeEMfiy2LH2nRrVsxTK5kvku0HtfmiNdDr
O3B3RbKWz187GyVVgKIAB5mXTK4P3RDMXoaRQgQLflbcWxMiKtUetY9/L6ioK2Z7ZuJl5cbjYLyr
PxbBIv3p5JZGHzOztTTg6Hdc6hdQDIO4qq2VGCMZJegpB2+UdZrktUNe0msnY+qDB8qgkqBRoA+H
tWm+30Siz3hB78uiQvvim77s+Yt4keWNIqIqtbGP1bsm/XzYXoMuWfqZcv26RxHODIHqlQmF/cbf
owmlnn+KGjyduexAQGIm559Yya71tp/Vd5mQ7M6JxyAtHscfXIuE4V/hgzyrXO1CY8QiB/Ue+EMb
LGV79UEwz1f8T0OSMizghxvpPovGZsvKu57FuJdzIPXWio0mTMKNQEgVLwCZo4Qo/qaigYBhNggU
+R8kf6Hvc4fhJCha1qu+F5ZDwTBS2LcI2iHicE/hS7Em25EPabDI2V6uEy9ewWjYtt1Kcf4pJdy0
9gH4+pZGw2GrbwIczy+5UbQi0I4AJau89W7RwwVSn1qbptFny/r58GrLgGfdk5d7H0fVBvNn+mTT
RWUtpmJNEh3UQNTND78iH/dLGyCrfV6ZHI+msOlROPTVcfdDGYIaBLyh10GxcjiARG2SANNYBFjP
wMkcy24cRXp1AlnSrLtwMc/06bMi/Dn+nz/BW9H2BS3GuCdMAejzbvSOHxmk6KA591McacMXMmpu
iuEnt/CShvSsXry5xKuzR0ePRP9+upd0cB5L0Xr2eAG+PXgjFYPKE6ntpBxUZ+fi3rEb7g4szb7M
6WtfiYyOZqs1lVNbeWm1Usz2qvLsBmivIZA22vIIAYvloszN3voFevlytYiVMO1I9Y69P/XRIPgx
wsr0Sni/FExkC8dVlkgLRVeFJDb4GlnG5WVmEdUF6AtfGf57uGBjkARIZsRRzUPy8L2hj5CgxbKU
cFq+ARo9JvKfsNNk/FkV+UzwEgFSoskGhcjrh7qBc4b6YlEBh360xjEyuYGabXLX7d7qEK6FLKeg
vWAl2cAmEYaMmqZBY5tI+aIm+OrGYDEuSqQJm9MHGe7nhfE3ByJQZx0vrmBOZjm94osZazVm8URU
7XtlduY1z7OXHUwf06gqNZlb0/Qjwt/BIoCmpcXjHlnXn3818PpcEOpuZTQeweTF6EBw5+8atKB+
Mb05WE2VNGeoWsSkpbSvRP4SU2Vuc7URZjDsBXqLjZ9FIqNs4+hIRDPViDzbVgTE93teXMBgUQQI
g5xDN3WheYjCjWFpnEO8kY/x3bW4cdbBFMFho+r4pBFfOyzx414hQivMqJwxBJprCmkJUPKcENfn
prNwzqTMRVLOHVMISjNOTpxurdD5WQTriS2t0qW0ywWu2fV1CTBSa4PCvL4++hUJ7SMuRMZ7VmSq
xwVNXh32J4zJ6JwHYQ0bRU5sVnuBS6Rqod1Iwze6Zwe4Uem5ZU7WC/hjXNpAITpuOg2lw2ak4JXT
QsE6qsCSE2ZeO9u4j0K8FuNSWT+WN09D1GSUVHOEou8G4jdaR1CJ+ClQQHG3tboA5k3xtJ18UZFr
CzRrlk4FmrDwVwfRmKHWp4sLgNNcWOTFVPY+Sn5RxHOrXk4nE9BQDyKfCOw3P9XQJ6nyaS/Iugze
qg+GGNut1wirMoa9pTtRY2d3jeUgCRKgy2zX29MFOy2oB84ukKIMWJGJ/HB+2jbHbw9dBluBQcJX
N88nwaPeNbG07BwEEy3O7lh6/pp2zpDfVYXfiydl4tKdI9uvQvh8gxczdBfBqr033hZZN0kECD/X
GT1SutY4nzrh4iS5kkSRAot1WsGnELLS+NW1Jbl714C5GI8oEipCkIq7Dbj+uPdSr/wVtnqzOD2g
5FFP8Zp8Oq/TYV0urOHjUVe1uoha1Os8JbxjDMHZXZmAfkHRIUooVbxAxxRCRokKZtHAUpYc+RPv
OTlolyTQRybVKWsZ5zLK3KEGzn9oRVDLbdm4oozfyh8wOrIP0WdPWzodIabokovM9KYqMqI/JgKu
XEApxZilU4j6SY5bpuU1h8aBuhz1MAapSK1rJwoFY81o6ZDuW4OpAvcurGbJmOdzohxJMYqOm3UZ
rBP2/7kwna521EVTjTp08frfJ8kriUXp8gShu1bP8+v4BYi9LRsPEE2+ox13dif8unaUs0sm1Y7c
+TzF5kTQqG9SVk8qrX2+hnMe1zC1Mt6MNNVALvP/Ly2XnPKmg5iXdvaQB1p7fIPjZ10HNGwzcb7C
OCtm7DlAE56I8LZERN77oTk66VWUwZcsijdT/y/Bp84g+mBcpqVl1GZcd+HaUDdwx6bSQ9IIMFMF
V7l61jbXSTu1iz5aJuJxNJU3LpHeik43yIHFP3Q8fvos5Nz2ZXzWjTyuxrZOEat6VtF3y1lYWy+H
hhCeyG3C51vHK8iTZuChM6R7o+yRlqyE12wRYWuFqwsVw/2yXyLtyFhxJ1aaezsuNFDIbANO98Ij
mAhw/v6Ho8zLvRXuN8VaMImG+sov3C8r/Rou1bsCPneT75nkTaFPYK2dXlAHihYtoFsM1NVO2Wah
lNUXhaFdoWXvqsO8idGwHZ25NOs21bWkCqtLFL8+zS+r6yc/VOIZ+xXWViz2ex7gNwknc+ZM+wHO
Yg3DU/hUbL4YjGVdPNrt0/oGxJtqextYP2Kz2D3sIBXQPt0vr5iDMGWKmbcgRRuMDkKIgbqzK9qR
PQESNl3UQvfpvSzhiN2rVgXg4ZTgZnMcqQrILa8JPcKTShW4v+/6QiPBJo8EIk5oSSG/n71LszaB
Xx1/AlGsI5eZQRzBnMIz3TUqMR3e8q+vo1vEyg+TGjNNxk2Pqyyq33h9bCdApvlzzjW7RtYz8Xnh
yOl3CAEnnXOPalgqsGWj+weKHUbG5nCPds7RsslwT+0Gwbmrf7RoAy2oIebni0sX5GAxaMO/vgxR
MlemlMMpc9u76S1ZbgCIiWioBk1p24+IbnZ7VEkQuWo9Un5y+4c/ETlZX3Vzn+crx7xAitplBVcy
I8pnJUM0bDnucLa78ZUBurHcoM4A8EbFrZLp1bdGHqz1KXtcx7Q5cRY6dtXbmk+jDbPTZX/Scvq8
hqdM8uFamsqh5nYVStGsrYcJVWi5boetbUr07hUnJ4oY2PMVrt84X0oZM8BieXrlFpql5fgyfciR
hFpBalDAAr3FNrEew0CkU/jIymIpn4MH9Jppbxc895yqzhoQpsR+BUnmC7j2atshR/GGcooRp4Uj
3ndKBFiG4coK0Fbl/Zv4E5T9V0uuADA1f9XHHIRqB/3y7pBFetZglsZZLeucLT//bweDbY2k6OTe
ICkI/MrDtuEap1eMMrtitvH/BtQriv/iwtvvDhqqwl4bamzeZWzg8YXgoC5s+oG0lN+3rvmfGL7d
+ohapM/So/J/OqbqGHATKhq1i4CIf7V342055XZRhQ8Pr5L/cEwDXoR2dIHV3L08LaePK+IA1OZq
MxJz2ljFr/OeFmwXRcL6h/+bg4yF/TzJ84CiMZ4oxcAzUlwTg/EaWVVM/j6xIQjEm8zDjKnJ/YZL
eeT51W1XdMF7aWiILlxOR6CIuKfFhF/tnOd1KbsmyhnwS3c8z3n60heIwQQc0EWvixRxNspWDwe/
F0ytGcefAVyY5JV9dXUOVZUZu23CA7QJE/HR8MNWjEOfrynNFVjDBXkgzBL3Vmdwn/iEW0jTQSb6
RTerIyJEmg21Z8sPLCy+jR9nJWSX+aMTnYmoMnY8SD6f6dfVaFMI95agX0VBHy8ANjSAlaWGTSOe
h2CE/En9PB6HfXHtZ1/GdLEba1K5T17omHWn+L4hlUrttXc8sLRDP9umDcI2i4GCjLdCWT9y3Ptd
roeOFV3O5V9BOdym/Fu9iLVJN8BSacOn+ClZoR5dBC3BO9wa5V52Fn0Vs6tuYs8E0/laKqv3MLzS
Exs6iMkSoHKCXlIeZjqj8JvNbymKrOUZI8uabz12lcAB0iaMF3RxUFse819p5YqQpT6e7rw9skot
E12KsI3HAFN2urSlqq0SIFMCfrYkJaUDTaSASjK5N8/H82Z7D/s/WSEisfGdWA2ne0Qa5rnn/EQm
CMBXbVgRt/Jj+Z4GovYx2z4+b/6SkF9wa1/haAS3VbNUxYuF6chqQ9Be/ewW69/0WYFnP5xx57Uc
38sn3Acnn4jtUmWpEDc+GWdAkloWzCxk4YPPGAbxooC4BEJZ8GbKV3Jet1cUIY4f25hIlRp4tjA7
st2yb6LkFB7R7YwBXaovp4pOcqTPShLMd0sUqGdvp8dgVL0QI7AP+odvueknJC+BRNPUfXF1HOtI
OBYwq+so/EVcSUEs1Y6qx/njlYIm9f3BEx5RO0BqxjqtRdaARkzfKvZFRb8Y8w4JSr4Jf0YdaMiu
VRJarnYgliLfwJmsOp5FN2Dq8mR689I+VXuejoJ/6ADHaNQ3kEj5Z7iFm3UpLONlH3FUPwzb0vjS
Rfw7GJxvSmuqwneEBdiDo0clH7L7vmeThWVY1Z4eWpS73AnqBJeKIB4MVOahrqFKLhCYUCStl7Uc
cTVb+uJ5DRjnRvNiIf26HCGFCX7NR/cA9Mlb71VT1g3VVVX3LrSVUEsNS6holmd+h4O4xrtMwZo7
1N9NFxgrsk5ZXq12YefPFrZ2vtiCmEK6qMhSn2I8OPw+7ttEATiYrZdHk98qyd10UFQKhe8PayZk
WohBpYF+sA2fgWgO6WXooP64yuR7lfYsxbODjl7YP5g8BwNmFnL0iFsjtRyBvEOmZ94EBEMe+58V
U3xAyQkDGdMV28KfhElyL562+UTVJjRfz8e9EgqHIRaL1UBzxvr0X1rJwmDWZtkUl84uUij+EJCb
gqVogVcMRVYjcG4nkNgBFzJERYD9qcrMJ3onaNfO2PPnt5aFwPuNYvxztQ0x4Cf+f20W/lDHZZgS
Tm5jmfYt3zwVtYIYjADEulLrqAy0totqSINF7XbDIzarPuNF+vC/SJinGUc3Q52u+rJRj5vcjAic
W8oLLaiAZ8iaxgQ/6NTzLHqlu8XOpBXNjf6YXtwjGjo+Rx3mMnLww7+aqO+00l1xdAlJs6pFuBXc
j4EGvZxvCZGGu9dI0Md7fW4plW+iQQ0t3OnScIzQybKke1IoNREMD6L4tsgFb1fE9o1l3RZ68xyc
sf16HEyNA+V4CS2SthSXbrODh/Fr/0yZqoSkX3StWzMoMgm/SuuWDMZ36uLEt9L4XwZsYkp6LMYe
tbIyukro1PE/X/LCJCC9cW9YZBBUrWWhAxxzRnxLiTM2YMC9Zu7nuof4duIHHFbC/irVt+duNrs6
03g5yVo6Mg3XJ1978yhueX4mPFV5kzMYFS/PaNAdXgJ5ANHpBiDdkCDNbZZ4m0+vb0bM/dFF3BRS
h1C2GBuxwgJLwpnDaOOQyrXFHkWniWvU5lilPxbkklZTEsi7cIrYGL+L9w2soqX9bXG686hdjI1j
RtEsG5SuyXkG+/eRY2BhE/MNg02gwzy7BcjzCHTvh4oHTNIjkFXkCkaL/id1OydPG4VpCk6W8K8C
qI2qZJiaK0KccJKqm0bIsPTmxT8jHX+8D2fwn0RecJtc6ZlTyFF+tkPgmsjnW8kiQOraPCSyHvgH
fzhn9NJ52JK7HE+Sxnc5HepNfVUm4jcGvjhCfpnDMeTL0Lg8jOValq7EkRFnvfU3kYw88x3oZmvR
S3wCWHoMzzGOBOeky+0MTrTiiFxO3fyzPjE/LZy1skTpq+9eTNKguhYTUTRBfWkND/9azL+MiFOJ
jENnfbMm4zcf2AYW6n5WM/YCcdE1cK3q8fU3XcBG4N6CnXDtZGKYNUn3G6jsGXzXJQyWsXJrOo/F
GTRtfnoNdM9iWBzUUTlosVHBuEIEV4eirYy9fvplCwbzDtECxgHpKMbLN2IjwQUDCuq1STxTwEgt
k/enV1xHVU8h/cdR0r4S6TjF6uMXC2990WLvsi7V5AHwdwL2/VHi9yjXtTlsDdR8Omsnl/CE6Y3q
lC+rdfoCuMvYkJ80ilUlX7VLQZP5ZqWyx+cPO57JlwD62jH7qxBgFroDpkqAc1sbLRntE/U0l86l
OZUbnagOzSZngoImfe9rAUNVpL4fAVUfxQZbWGVHzMSIAV5X6y0RJGMc8h+sJDA/gog2Z9LEG7S2
Eo02SrZ7DqBr+95D3ZImkZ/tn0NhVAhhOxjgWzGiyz8aW4J4DuLEdQ2HBP1zb9wFm6euSqr/RDPB
27bJxbyo6IFpeUcrap4ULlLbvJFrTHqV11NwMP4BZtKQPr9Z+6UbKwI0j8Oc2eLxjqjhqh1IA6tC
OTPTvARoD8a3lmEIRso+WM4wrpgbHpW+VP7yV+FO9vz18hCWgURt5BcGESCgOPw4KJUlg04iA7cV
4pLCibxa9b+eF4+e+WO3VLF9cJJ/5SAz6glsYoEceMB8mEK3QR13lV8X0xBW6eZLFR3NbDtKxV28
C6QRcMKXfUq5buy3u1/6VxusHkBHnaRRZx1vriQAwpCCFmqGtNaiy3eoIAvu8XY8xuQ8JrqnrZlW
M6CoBhpViozc/NglcApc2mFFsF50wquUw+Gj9afW0NatG1pbwYvKzIr28ryfevyyGbT2/R74ceNW
FW3iOu8cURrQY3Excvb2Fv199swpX6eEr5phchOlryomPGv/5DpFyAba18YsKaASedFL0ss7o2xv
qxazP+8xFiKIPmPZmZ6QWHrr4uZNaYTV7NykfgxL1RJm5RxYnLCD+7VoSNwKHoyZES3ovST2qN3h
qQRoobis/SLkgMti1mu3KduXOdyb8Zi067zNFlr0GxG+M2agWp8cf88dx1R0AE+G4sj4wI7eUFFi
qXMpKPNhACUnNK/upQeUEPuTogxGhKsoNm0jlAh5sGwTdBxZCcaVkZ6brb+65sc6EzR9p8qGpMCE
WnaFsUeJPUrL/COXZOVOIWakkzIHZz0L9deUbydMew/9iPqGPYTjoF/SrLONB35Ldq3MbsQ2lHGS
IMl0k22vtz6HZ1UdIVel9uupB21yDQE5TDfHntb7uTD+gxj1PEybSWveyGSnOZZMr4AmiYiZCbol
iuYCSTNQiqcBTiPazuj0vtIvZrO949Pbl7t1sPW1uZEbIhV3RNyg6/lyt/eOjEAqX8V/B/Bqa/a1
MhvZLCNT4Go4fcO27bhvdt/y1CBdN57GiZmBSKjG8W5UTZ9/hwnB5NmqZNPJrY6cayL2O5ZnjjSB
f5JYvHo7t25kwa3G/q3OEEMNYeqQz9IaaXisFLDVLdyP74GdmXzC0DcqOJTNXM3zW2QKD7FTZayu
+M9alUgZtyPBgVeeaXgxA7q67RLRmSENebmreOix5zwnl7XEPGV1/9OmMKsoEwgOiKhX3QWhaoCe
DRmYNCrJuk89U5oNWRCuc/aTRc5emhaKIqOevomvtax0zjpT0V0bcAXlVL2FOKx8GqPfTHrdhFx6
yPeMJGbP1CV83vDD+zOTQJSfsU0DA7J0vGTXAWz5D8560Np39cERasRh44MsXbi5Tjocdkae+96R
7XDl87ErdjeLxbkkS481VhwSXoyHqLRCEZFinq6bBXf/tGkPZ605pjD7ysR9l/v4J6gJCOkj1U4H
ZylMKugAzncUWMu7HsoaKef20qTvhzdK5X5WlyivvY1UtIuMNdnKaqDSBBlysq6pSSX9F2uz5x1+
QJD0IDi//VbQ9f+DSIfUElKtlsu4NxJK5h3SA5lXCnC8RhSmARL3T7MGmLTsHZozYGTtfNvNHuML
Mb34lOICmArmnnTubBkkIwKerEefZCiOlBhdxnVNC8jNkHpbVsj4Ii3cHh+AeGE8QjvZJTU4s2E1
B0OLAZa0kt/Vp82KnFQOHxk1H1YaejgB5QbxeWDPwVhfoGnnnLggQvaL1LbCzRaDQp2aAzL0kpQp
iViU6gJV3I0TEdM7BfqN9McnFibnfDDr18XF8IIBscLKxCk87uiryaVw4lYr1jArFZ8bN4YkWANp
ZDApeOvW5gkcoluM+ZSYcZJkJ0yfkW+ratav62adH0qkRh4KOfHgJ1B17zJgvmnNP4TiJ7jonRqM
BzBh2/jtsQ7XL+2O4tD3QLAjzF+ujM3QLXxH3u++2CtirrGsLXZRmRLQLtFnIai8ReSYFrN3kaoK
mTnMW/k1VL9VkoW1cszhVVFlG56yTFX8yUSo5ULoXf7So3Qt667LP6WzPAcYTOoRIEzPT9Lvt3ha
kw5hUBVhXhGgdk1Sv56EkWrkfQqWkbFVscBwN3qFBIdyqsWB6CNfGiNj/5qtsIQKOEdPqPRHl2Wd
zEdAwzkeJdSGFV7ls4XgHXsHY/sgOWqLNZpuShRlHfHXahgRsV+s3QhoOiKqMcJqYkWrIkhrDtR1
sE2/zOlXx2nqclEPZsemCFppemq72lvRmqbDNXT6J2OvgMgPxro9/KSCKt9lL7xhNMZZ4P/6eg6f
Q+SJkcndqlLAxLJXs3pskD+NRfcUWopUUqRMoVJNUXkrK1BLySZy6QL2LRAWuqpkBFsxkeaHN5qR
aopJRgF4C/ulxjGG4WOPidkqQ8Kn7IhHdiQRF7tpZInPBDczo9rB39ZVaWh/XXHml/1uf0rKJ9hp
XpvpbYhxHkoh/elTp66YlJLic2ibWAnOGG4EJ6C+COWtHOT0Se9vJw2A3ua0wmtCQSApgSJV4yW8
fu6k1XetKPc/AETIVDtdEP56p2LO+kyoDq63InxxIIwbZTfFlXcaqOvQD/vKWVrNHySfVJvlajXW
oI7U1VOxLHWxPoMut6V0aIiAi3Fr4e/eShDbVEkJ4PbOngQEFOGgrdlIKj6JgIxrAfZRONBu4j3l
uCXifsxW9UxGu3sFkuvLFYBmAdCMTYZ8KlH71YNaLaYFBrZ3s51qF8DBt+xULJCwcQX9aRgurbKY
gId/nv9ShMnvKj6QeU6FzDUAAHOh4Ac6wSb9xhcUNCcIm6Amt2F51iFEBH5A06eULI5bHzmh5G/R
f7YQAygq9dfSpqHIk+OhPC6Q1S8n2aorZ+1lxyvOXg7zOMKXcg/SDUo0QHGmQifc+xxiUQiFrqlp
U4qze5kPXVkhR2Et11d3QD9CNYeLy/89ZeQEtgswtDKceRSYDHbuZPt099eC7cz2ZFetFlzrEFGF
PxB34cbMGjGRNC1o4Hd+g/51/ywdXOyYjlJ8mZ2IuYsF1LQV+33nJS+dxpOC28d56Ho1bWI2zjcA
ETTHRmVT0I3+MKulNFlokxOgDprYF2TjDONBIyWz+uwaKmBuoTCDKV5j9Cstfe0s/EEcXRjIDUnn
4AWSLQPVk0pbQ9GBVlE2ol5ht6EAcjuoHodpXKS32PEuHvEB02gpYWeoFoMiLtW8irWQB2bmCDj3
Oy++Y1jrt10A0RsGUVmwpys6VkQgblFgZ55K2MiHsx+GjbyDYcqVbPtOWQwkGjZgbxk7Xx1fLtaC
Q709PXta6kyNX9Jr23UKfwOXmztpy681XN+Rclt2qV913p3aQ1NK+boZLYAl9zub8wH4fTMiUV1C
UphfYtUSJPOmM4fCRgO3kPXltpXRjHYbzPdlXR3LfFjETHEweezP0OQB26dlhE0q6wbcEXrbyCJr
5JHEbR8iylwlHtwIC79O5Gu1a788tbI7D147hO+TflmCeKaUp7utZDztN+CQiywMbJG2IeZdaQZU
6P6v3VBtThh3SbASCewhQG36DE1SR92X2yLnLgZmtsaF66MugkxPVOF4R0dBSNEgigmyh5LPw12m
8JX4/iNVIuaUVA4RpTQ+I39GqwiZllzZoIwjjtp/jH2KKMCJGRemb4MErIRxMFcWGT5zs2meXvds
TbRRkensuG9m8F43AmGULZu0Dz6fy8zpRRj2WemZBfh9BVSsz05E1/B5tJ4nkqJ80hjtw6CEueQe
LvcYVuC+DUWyjfWPp/Js/SR4YdIsYlhWJKjl3gP/RU2+QjbJMs2EohYKYnQ7nuRmvL1GU9p4OAZ/
yaczhIxKljQpiXFRMggisfEr4dGdHCeNrXs1Vim/rSJl7qPYfwcrTtc+aW0SDcQoLEZPdJ4SZX/+
QQIO6PA521kvaOm3s47tvG4DxN7f10fDvKFesZEnAuWx/F6NGFteSPoLH3ajPFwh58eYmWcB7LHJ
vGmj+lJXg0ygTFIHIeTStgh61gSO0+QZgnC/t6lXdrSnpkKqvMRnRz/Cq0OS2o9egJsGIjw1pSYC
tHKjiyesHI4+8NrUGEI5miK93saYIZQI1A4bf/hdcWxBQflXy44E2XBbdzvjKf5SyKDbrhu6tKMe
0Zli/++fyZOO8hr7D9v6igq2f4geGRDoinJKPPNE9PkiHBQ31ckq2OhvrPlKcK3164b1eS9n2XxH
TJ2OQEd1HDasMLhyArf8+AZNU72ilnN/jCfPxwYHkkuxzSxHU3FuH1kY3zBPnMTNETga4VYetXXL
h8Xl35trhfI3hwyIzCvBmqqtJFJ6Slm5JjrCFFaoGZ1ZXa7Df/jLtzLsw9mXkT9rUAKxCe7LI1vH
F0MoiDLR9WMFCD2X0J5UwP+PfiklId8rqv235qZ5V87dTeTXK1DxnbD59Y4nrQ1eHq5eR3GYEAQ7
IXikvJ1sGNFLDfO9/5FePeeXP8nxMqzyUcJtDs+u2wEPi+p+QYZa2/TqRBz4XwThoYwPGcMDGhxc
BgLtYdY5q+ZNNdhF5q0UEqQxtICg4FaJFLxGIUk2O0FLD8iTJTu6XgDB+NNxJr+G3hV8RdxKaOfB
duRPbL0NlN+d+h7TTPvYOTigak0ixVxOVER64TGItzPIIFkYLsgO5bFwSskBeDKWxxxdIXki0sBn
6PZ9+AGMia1wwsCufPaowT6kaF/UEMMRulljfBeA4ReatLBfSgIessn2Pg0MBkZlNGJalYhu6UMD
UUTxWohjYjJ0ZAYsplKNo4V5h5TJlDOpMxGH8xfsAB4zmUzBIxOGhdjxqGaE0IKjDqKjR5Zl7G2u
bT9ZFrRoyWNM/yJNfSOyLllhCVP/QLtSIKkNI6IY/HZvK6W6LfceOTtgiL/A9v3ANHEZ/016ZWo0
RjFki526euKn36URWEVSxVyAzOZbMzc9QO4pMvpuyFoNNQaj4NhuOQ/06MBPc8cLXRahiH/9kClX
Sr0HaYNcN2NxTcZtBXbWoydSANdTcKENuqUsc1saCDLZhDjiD7002K9R5iGNFZRFJLr5FHksGh6F
boAeFXzLsb/sdy2fhMUxs9hula55kXSMQpVE3zmFYXTc8HA2dQb1wGWqjRj+ussgyFUxcEz0DPS8
TCO3NBlivzZtyjqFhrO9lXaTKTwYWCWZ8ZulSKClt6HsOqUzVqFMhUnU40MKCUtYBkRyjTrcdSko
OnM7GdZlAsIq7+/b0SDBy8hvjlYro5wulLyY3iQlbwjcWlBl1txL6LBDnJpR8U0bXOOM1iP/JfaJ
bcAz/Yq0r4mpP4wQLbQvwF2lgbfNUNPJARItx+lkU/cM8GbtvagU1nQ1Rhg/UtUYwOZdCoyJGDHB
pqF7gUlqrRcZAxi/lT7IKEIE4x7l+9AqguZz3gaNte5CKV5eZYuHm5JOQlkteZFEflXrc7lmaxVB
dO75Ostms6eHs9LWBxOtCzSeXd4wgT7uTB08bKkfuGYqv52rtF9WkHgjZN9AP4aulb1BEqOhxhNm
NIAvdI+kd9x5+3sbqNKkQVOaCOY4jKNtDVAQsOeASJ7pKNRA9Mm8G7cKha8ig9eQA3McXaBYO0Fm
osdOXn/YNQf0vr6i5EPauirLMuKhKA79M0bvviIZwqiX+XrdEOV9sbUdbiMBAZwcfb5vOgKGtd/6
WO37eObJvTTlRBFv/zw6k+yM9/PpMK33PngMJeSN7tp+qvT8HVaJRTDEkzQSBuSYhDsZg1HCON97
+nY5fgIIPr4PAFoVJFul2ksG7b623ov3Lm0/9tAFKQfxIxH8yPW9Y1ARmvCcoGmKY0TlfQ5NUoTZ
nomreklofky3COZzrPQWWUoNDV7p+yzpeNgvT2CfxhapG/YFUAmvGSPfNKrzaHsSi4+3RchHTYzC
VKcY6scUD+dwW7NcnZllzPoqh92Trso+JT1ZnEYf4mRSqkeIRynJuYTgjqjFYUfVBGPMUC4KVUW0
O/EYLlJ+KtKUK8gizCNUhmjbfwqUDtllEmI2jJ7lE14lTZc3rEY6q6M7ndRX0cjRYxBSDRwDUpB/
MPPc1YjudgWoF93zVuSl3brTF4afu/kHO5uc0EE4q3tCA0+QdBo5KFPyHjUx7SJWmE90lSIwmXjE
IGnCwKhAfeSarP8RwJHJ30McaKYagq8sMpJ+C/dtSNmf7ZWco60KOtew3VjtF86uUNer6yvPowzW
zJwOGc9H+ib5mVH0iKQhY+ZNLGZYWEz2edGVQFN8e+on+PD/g3rCV7j/g0ABkWNhoNvNHxDDt7Ah
SyULJjEzhvlRTcYTNRnEEcZGo5341XQdqzKoYol9PjKHApcEZ4A+zWo4FbT9vZNkcs8qWEssVvV+
hahOEb0JLzsuZQXzY7PwjPx4UQXxlxE5GyUfIfMZB7ZuqZ2G67O/GCkY2QO75BChkTApVF4EPUtK
WPfX7evCyhTm87QJXUutIKNFXujEUelFwl62abPvSeaqQHNoZvPHg5EsxGFEnWKbD6afWbtVRuDg
a/D6rMWUujWsC8FpUkAD2+wIX6m6Cw6zo3WAYZcVKGwmGcI1mGGrbBlTXexIEaJz3KTgOZYma5oQ
dRXp9vTWronLuLSPOdsE3dJNjXR4hrx6MAiZWxcbkpS4TMPv7DWw3VaMYXNv67U2BmOiLHZfJ6/b
EtZBBNZX2Z3b/xN8Oo+kZNSSuEP6+3OdUK88Xy4p4wwA8pUo5jSmdhTRh1VEFsi7RprbQ696YLFo
kch3pCiHa+pdWUQeiWe3N+7ZIobiKzdshk5TY+8uZDsepnBpQa1gOuct831WLHz2auh9/XJDcyqJ
MwlRhisftpqI0KQSpT9jZa7/VWrqhSs+G2pfL6noNJJoBZaHFKEDgff9/3aCasx7jdBFQ2cv2eaP
9GMwrg8Stxy7l4t2hMx/R9IZhu5UoEe0Nk4crysUXEb8pwQOBTtHa3CaT2e9CftKXsekrI/MveFc
mA2GIaJZLm33bXMWIt6DgNPS3Bs/79rK3hvQ/s37wkVrirV95D1G4R7YZMNoGGxCgbSDfyHwr1oe
AdBj4V6gBBJQx5m5zQfta+I+1OzSEdisnd6KZjanwQ4Sn/ejMoVsrrkQ6356BVnBUukna6c8VQL1
15PiCkonR4fln+2XAtHESjwazWvawn0ohfvVQPaIvfE61Y9ZxHYl+qIfjH+vjAAn8iZwwNSD0zwI
ekdfO7VO27Y4RtjInOlS3aAJ4WQRZtBmof04pwPPh99+tUXLj7rq2mhD0m5o3psP3+QSaWryLlO8
ZmkNH8h2fZ8uoPID0NaVJB5jzrZHnws2ZbjsTVq4EtLp91Ito5+ad62uOTQCKFMIlrF11PcoW14a
29xovJKgUb5LGFA8uC/zqGr4+8U9M+9ZwYj/LVzyKsHnZxCPXGWdwKgWwwv40zlGfFjITKCkCFL0
A4qTwijQySD2qAvTQEzRpEEyAQaCeWug1b0xqJRKOdMw7tCORhfDlVDBqUo8YnhT87Jb8gqG3Mnn
AM2xmeS78sOhYjVp483KOSHNMc1DrIx9Pe4iFkDjsf3K0PZl8825xach3UnA5O4bl/nOdN6nx94P
w+ygh/cSzb1jq6CW/n1HD4MHU/gJ/63WGvGF7UoOeW8VY6TGbmbI2w7b094AGDBZAbxakmGFO1Nl
L3k8tVPzLuinPdpCnc7YOpZEvTocjIPh+DPSTc7Yj42dHIWEfUkl1khAdxXRgykWPyJcbbeZ2YWD
nuPwQpWFT6T3y6E5ave1XmQy/E12EBSH/4qFIrjSH76hgVboi0gglA+F7eKF5JYqNjqqt/fO+nfN
WaOqxs9RTLS3t18de1sU0ragm5jIKJW+1zjKqu9o9g6QijhnYnIrN7xI9dQokggSx3KlE+hsiGDQ
wWFPkF01qvcf7psHqJgdNganXP3OerkE+YX2pxHdjxKs447Z00mLTlEaCvZ2wwFtkRXPoHNAEzWW
or4HTrM+cltTbZCqgU+erqz+kxUyb5O5rfcVKGsXvBhLHlPFxGWe6lSa3AJk+Djl3fjs387pP7D7
SGwkSRvU0osr6vvVy5epnXHH4AMw67VrJDJxuY7v/Nzjb4uHq81Y3E17olqpetQPSGoS8xTptcF4
L6wx5KsKAiZKWOZbtK/+i1Q9yaA1zwsnBMttk46s4c1VvvcqVo9MmISFiSVPV1dYXJwyVCN0chsz
pkL2jEZUutJWzywFgsxYJtKg3PCRWLb7SrKtD+a7RiyWnRBMxbHFRXzufC/r+PVH8j2TpxyWgCcO
cKYPmtPniU2Sv0l6EJsSgwaccMptzwE3GRI9W/aG2zdZCfQrexW1jHjzjFGmmbK1nrXFAdOBO837
epVrM/2n8KuaaaFUGbdpDfxw36mxuyhs8PLBG21fwyVLA5KpTZWt7+FtBZaT2TcgPpWM1AqPy3ir
ZoCQ0LK+zQYT9PE/MBzSF1xn5gpfuQ4hb9rcHpr0xyKo5ulAbJs/tzmDZCxIt6SwMBfpLldOhCmM
Joq+WNMnJ2yMr8G0hzqdGDMU5Hm5+Kn+p7A5TZovG4V7GkIYEU6aZcBplTepZf3jtkoZ+xK+sRpy
/76dSmSAVJ/oyy/0z98kthlFXggt/G12y7z7IapW49z0PxUStrawKRfYsjuutdtjNP5LAnGA2tK2
aJTKV90BP9x3dbCyO2Yjq+GgRATvTjoCzjTXdC49f+gHBLQcGUjaFb1yH6gLVparXq7XfrDXTO+z
pmHxov8HqZcYtyFiTDThVKI6Yf2mzkH6hj0YxUUthMCwuUgqhhn4ZAAyDyyTuIJGsCRjZH1njrye
3BGFC44IMkWlF/UcwvBwzqwmBvxbYNDoPdRt5zUI4q7dsA4LMH2jiGEESLuCz6vfjNXaiT19SLyp
MA7Bb3dJyLExt99mOlILzzsjkiQbHvMCBDCyMK2SXEFmMuvb0XKl/LCPSJyHk6nk4zE4bAx78SoI
VGTJU+GTn2X2NNVEohA7c9lMSHGVo0IicodGf5XUNyb5KSJwwuXJ92NlxRObq1aWrc5xkCKfVKf5
86FFkQuoCAWkdGNWqecXJlx/k1lnqzBlzRR7hDu0vW37Af03isRnN+YqUtROQRiWL5XBZdiqCfxM
QfEJYzZY2J2QvW0gcam13TAeQWb3v5NR9zDW7HcXbIcoM62rALmqx5y47gtnteOpC0navlDXgBvG
NknjSNp3BKvHsfstGVSmNq5boj3vfUgoyZLUAgtx2ye85r/TsMuosAInPTjyO80ONg7pfnz4Ts6g
YpQ0Zczzoe+WIEcvrzk1MBEd4S0jy6DNKH/03EDMwaiMbojmaqZZFUdz8PHO1Jev+P9MT8Hhk5oH
Hp4DSVDNYgElUXJtF6AWCy4En87OBny7uhEUgUY+w00m63zcnGcPzYtwdSURuGfyl4bM+zz3WJn0
HWMhIYzy6rOVSenZMtTBQ6808saw5TGim70dCgJh5KjFaSB9v3efgtsSIEMOLZXZ878QkWe5N+Dv
+RqfX6V4y35ZPao/x7EpeWM7PLVZqcSvbX3EgwsVy2+rsrK4IkyQIM03yBwTFqEOE6IVPiqBHycn
1jIFVCDLyzvgwHgLh/6xk18QLXG96cJ/mbjAO0tdNL8DT/eOxaTApA/z9TZ4d0nSf2RvDhJUeLzj
LXm6LIebT7LEbH4rg5Piabk9D/L5uPtwfJNI/32TqfPymmAuMiBwB38FEgvAtChjTymzb5dTwc4z
ZhVRmZWvMmM2j+FulI1wAAGygaHc1R/MP/zBUoslY5aZ/H3A88JjtTHGccnduR0Yhz0BAZg1IMK1
xYTuxIB5p1IyfvahQm5LDTXuoefGeYmLFBX+MsYkczK/CId4eziMHpzXkA8DdVFE3Zlw16+frlvF
kDoWYwrT4JW+NfLTy+gJrcCaRD0J/geCV7txtTiq4Y9h9gmzRrEZ8CG7uhju28Tm2Osu+qgrFQZY
hMiP4k6Y72djL6wWeUwuChcxK/rHcffOKT4u2ztwGVrY/7rhx2fYPEds/lx5MrSwlCUUFJ2uLqfZ
UQbJvZL8qB9oi+6Oy/i5H56P/1pfNKlIIlpoHFGhF6RPTU3jdbJ1Ts4nFSypISSPbC/Ct9/ru6sK
4SGLhiwUQItHvTrV64jqxlym1vLykfTRk4wX3Hs3rQi9zMOgdv1+f4KVu/3BWkQf2rHE9KTjEHie
SROo/J+TjQrlqqgQvr7r5MRuMDJnGRmKPYj2igfYURq5Xr2kAELiIJapY50jyPNC0qZie2wQJxbS
I1blWPCZXy7+CmQXRkjzxTC7G0o7RZw9HD4lcYLbKeEs8xnhLIj6GJEs9oiZlf+5BoPJbHC7pECr
WNcIqnOkh99JWMZ7ewvJ8WxZycfuCZDkujt+tln+rAx3DMT19sIFXDW7r8f3CVzjFSotSXOZtCJN
E2tA7fd9Z07rCUX7cA738769Rbr+bWfNZRDaGY84CPsHg1ZfzHu33Z6/O0DbuE67m0SZae6TWCRV
HMzDl2ayrwFmyllCbJxf/yuBo1RyW+WuUTFNvIkNvd3P7skRVi0VGbfhwOW5dwntQ4qsSmaLE94Q
oaZYYzi2eS/JY6hI5nma3RVv+vyYF2PbI+fmRy1rCHjhhaKoovmpE19Rf++M7U85ipxtOvsIz5uT
oRogohiH8mBGvbwkLOFGSa1oJ35VODw4WlYlZdseQTLOpVFDv9abmy8CAYcaJ0Kk/ugQgHs92S+E
iE3seT8riX3fofkW9SjFzm/sHCD6gk+QIBMCFiNoqq/YVrF79FlgylXxIhViUz7UQr31EJLiqLLT
Bwq3cUEInb3ke4L6qcXhpb1fJn8sa9wOiH0egJz53IV9OnCIr7LLrXIekzaShhCmYQFgvDaX+GfU
4olCKOvwIxSKeHnpm3n+5vOLzRu7mw9GvZgFRe3429IRIZempgAkbSYuoma5zhCyaghLWRt6hvOP
jkdNnDZVFDEtIN9Cxg4o7PTOZTqGpPDzZtFoFyfC7TGkkzsUgT4rY2won64tM3xhNj4uUKHb0Omg
IrFSo58En5mBldotTKZfbjys/4/jF7uKpyxB4yrv0rKNWPQ4UCKz7Nq5mumeY1XiByn9NUnhmZNo
VOoVs2gWIqRk4TKlTnlgYXyogJxZY7La60dXVcDldhKLQ/RV6KV1eHnHlopCuza12UU4uYm1hh42
AoCIQPZK0jfD+iRLxVIAoGOddEEcxhqLX9Va7pxvstUTv3mp9gRa3LQ1e2UV7G1P65Qnj9gsdFsM
ZAD2DFH759IzQMS1v82HiZt00wn06EWhP2nC5d0p4u0/xAmiMLlh4OSW7wlqOvDB2T//1vXfPqMR
xthGpmYNfSyTnSKJWEZlT4aOcNaPL1SC5pZVs7B94sSLnNPzMUL3gAGdtWHF+WBJM+LAAjEMo74U
JljXOUFa0YcWMeLVgQuXo98VU6n0J/Npq0BW6xN0wUTGnFH3BYfmfu8E+DzILKXoBARAFQhTWaTu
seIvz5LhBPQi3IAT6ME39oy4tgHK5Add0YlFhDfu+eQiIP8xwDeMSySWVF8Q17md2guXHmW37PT0
RnkFkxvndkRypArvF1dJru6kFw2r9V3Ts+78NfmM/lSpzlSZ23SPG9u4Rk/YfiGi3hDXh1WC6200
fmxd1rDRR5iqSWS5+K4gt0DXVWj/AoSTm+Lf7PDn8NolMGcYbmiw80WBCDDJg3phb2xh1hnuR++G
AI3eXqrUNj353G/DNVaJlg514pV1RPtZHo4vKfexShsARDhREn4sbc3xlJyk+p3sgJhmrnpqUUfJ
Rnqp3ciF/RS6KAXB03JWn/49NiqwcfrkFFfI7VULCDSUaMg+5fXiKyu3RpuHqcLrS8V1+uxXy2Pk
7vdjmHEatOtsxskB1ixyzbUIfOA6sW88iA9KeS32rWaVeq0ue8LSskIkY34HEtxeNifrD/8IAasb
p8vwJvvE5W+If3dAT7FBChDrQtiCXXv8o3+DYGlIEC8FK42sUnTzSIY9nxa2FQXm6D3JgPnlIqP3
9bw65Mm5Zr0YZqU6cB/h6+ZC0Sr30soI3+new2fnfhv03lVW/QbYq2vRVSMgZ8yq9Jyq4YZfxalT
LzaLc1OQg6V4g/hGGrMeHfgiTlI0YiqXPDg9ay5An/tUnM6Q5aNL9uWBRTt5ik5yv4ojslXX07kL
yImWqFn3It7AAbotfI33BWoXhId+RbPrWbPoX+/u+/8Og/qSiN7dwODjXSJSnrlJhnJdNKMkInzC
21xXurL//uAjijt7Ri8zt2KLhXfYFtr5B9DT0mPeCz3Mjvrvp362Gvy8ntvOQoXiKq7DEPGwjmRM
ICDkbVvQWsbUiyMGfN+NZfZVzZ0za1NMOWMAN7/5fo+fesb0naZFJ3+k+zRgrBRRUr16VePQJwzy
OlPHUABb6x2vti7RRAWE3YbcPV1KTRkiTyV2ELSKO43Ya9VBxevcKJKjEciBHhSniwNS0pqldBDw
DzHtNtumgWxRNGSAupPOfX/lC5UTlUrWQHRuzZK/nTjN05Zi5HYscL7cq2qKzyXdDYBn05MiHS15
47qWeBj9eDgG4YbvFj9Rr3aye05lI5C89FzM7qCVR8s+U2zy49Zvx5jzzaVhLvE7OkvJTyWdgXCD
MF7j+WuA+B4MtG7kEgaO446EYNY+icInZpW/eqzo1/lFyIa87E5q6yZfeY9SePMJHyoqq5jO+n0L
XTwRq4MPLTIQfWCPcArNqUoqT7wKkOvpXk0xJRW2sHqrl7487DEAdYhp3+YmLppep+pojlSV6Se+
79wHEiDl3BnhvORGkmFaNF0vYXIbrWa7qt4H2CulQqJ5UadKt20yjGnOEDBxgCAwepqy+e/fFwcz
IToIaULjArOK9FjoiosL/y64XrU2OFEm11fue3ef3M375zo8JHscBbozShV3dumg5GD0YzaNfDim
0gpoSjpHwS3y+o7lQUvrB7o37WJsVu1Jsa7uH6s4tS8kaahpZVpXKufzINMVEzUDmuy5kvYQRXu4
wXDMIvhJ/HGUteq72kIeGI6zJeea9AltzbMekAtPUJTJfDxFtD3SAHY5THDhqzqNCH72intetHXU
C/gqAXhcIMITlSpv2+Jv6TlDn8Psyhw/ldzD7Ho8WoVD4jyl4iEE1Txh1uOucg5lueHqVIsgpUvY
dnhTVCwo7ScqjcG/2VW4jCcR9D1HDDECYa4J2T7WUMuFoB9IaWlAFqbFrjZNKFQ6awwQmjS9YdSh
mzAZ9kgtER9dL+5PDtiieCCx9MNG1WbwxxiMKOv7+pHkH51OEqiaDaZmGKv4QnYFh5pKsGEYbEoA
8U1z/Gt8fbjTf8JWvvvdrl9eXOzG1MuxjNMkpDlJz5jycCSJa/0B9Ro3tknWwtHckOWl+6C28/ni
bQ4cuLHiWcl15rnOdbhsjLZDH2b3da338pX16TaGlgDjuhCmlzEKm8S8CTlRYY2SHhzarQD/BPIt
ItDBdvmNtAF+PXNQuCldEuyQY1P4DzNrTMUp5+/HHmB8ou0aCzWmR5Ry+YnJU3m0Hi6V7U9QLvsl
vyfvghPV0tCHk1QJBDQJpM9mk7edFGozKCEi34YRv1YXsxS3aHtPlhJk3/QYVhHsMNKqgX4oJLf/
/dVyzObk8nrF1tfswAq7bR1fIgtQnHkd0vQ124egg/hQY5O1Qb8P89iT+KTHYgALnKFM6UAMS7C8
q6w4Q2H7nUUEmWhM0EvV+EH2fAhEoXlkKa3yezvC7ITT15B1UOjy0Fv+odZLCldnqZ3176EdLDeZ
0Yvi7H1prgTihro8DqAPpv2gmceYvxAhTHW60jxcMfBe/YWS5gjc0m1RtWbqNlI9154huZchjZA8
DGCz1iX9W2RMJ6kOYM4doEmHQ+vh2ul0oGUHno2m57BkUupPH3yTgMyPAykOBhu0HGRR6vYur7r8
DqPXNq2qGNs3UTtG9t7PBgi7laZ3n/SfU5REuu1vMG/GptAJLC4lIE8og/5fSUJ9QYNRJWFXwxyl
j7UF3WPCtRkRocrGStTIVtS7zHXEDG+juePksX69xnajY6U4g0L3VtjoVliZX4Fg4bn/9Jk6qfKW
AmkvQJaa5vTsfIA22SpnVuhpK0WEHmZU151OD02hqA9pogKN+U1nfUeraJ09IMQmx7AhaR/sQVa6
1v25Q2sMA8VNHnHj9HSEKlQKdXGYUTEHQYs9buswf7gvK4CBuAni9Iat1XkOf5TC2Vai3sfP9iGN
m1lFLEiL+V61oIXzby375KKHDQnYsSTTquG1o+k7N/8d6E7l1SisC/1CSn0Xuiyk2cBIbIOWKnYT
Pq+Wnk/s6meC/2smAS1dm5fQtWoIsYT31TgL4J/EKRy4HWh4XLDiCDTYNT6CPAbjAIDIdQC6+aKp
7XSEqJqWQzOvSwm1n/0HzR3uZgNNaphgXcA46S7Q+nrZxpeUxauTOkeAf53arfhb0Aevxujr9VsG
63kIxDJoJUoSD6cBolFQEdvZ+tMxUKVyw6CNkPQuFAY8FU5SwqMhwTguBCGC/eGuXDJMb52WN/It
CBCKZrcspUPy6BFUnS5HQ34vMzVa0hvCc2WxUBPmevn+WP1UeLq8dsjyOLUJp9h1uddYHabsHI6L
vTifW6/kCZEXg/wbApBF7r/wbCk2ODdDdEOMVLSFRyKXPQqo2uhzyyLGJ7CE0mtgTZhmdK8LjBKW
YjkbN/fkRK55cQ5UUnCNv1/3Bgg9MdXCnXzAHkseDCaIpGdNEydTHOnVmqHQH5VXPI4CdfgY2wN/
vbBwjefPPgf/J+8cKwjgTkHVseO2TxcVNmH/4KByvV4WGjbxtTJ4c8pFYjU0hAV42bDq5XeU3py6
pvlX+VSBhM9ZgpqBM4qz6MbBo4BBaEL2Gm0rd0/9+ykoonvaLHh9ffU3y4QdqzovPbMZur5ApVRi
ZKUQT0NhuqSX11mvUmlMqNq/ntrQKbPrhQ1oiE+MfwSRPfSFW66zl7hmgQQHl4T6n8AXCOWVZmhn
9aAfRVMIpdjsKrSDQHn5r57fSh4v0rMFLSaSa0DUDrsOufKCNppan6GXQZCgGbk8tVCBGl6GdgNw
m24Tb6rOEfRTzUSDes+CkxIrjn2+nh5WmcQAj/cJPE1N1h8sSo5U+chJSB6yjt0n9KGKJ5/mGDrK
CrXU3gnGcLlAoRuCP5EGIfAOi00bebDohqScRKdcalfLg96QUj0yVkVdDbX2Ryij0EaWDxcT5FbA
9Xs7PfBCAbPbevbUSrtgJGjcWiVUK55XiWYQmxVskmGerbd/EnYyYVG7zpambWJk6wFccFpqwn+X
IpaVzT2pE0yKGnjssK45zmPQzxEanT7PLQM+ED2dWA17Y0JTwEiMuIHltZXFNQImEJ5P4ZRTyyn3
PH/MSJ+LhD68pMxCKoQ2F+gv1Lt0FliM6sSpbpK/RX1wd7tGS5W9Q1ocBAmgigvuyJ/AwsYdj6TW
BrzbEsiN55qdMgFHR1UwXPpvLlhQwwjwoseefwen50t3m404e6W3jtv3hVjWriPcfkrhmx68Urfu
TCiMKGktrI4JFwKdV8Z+sC5WRZ6x+a7zHXmnhqUxPATS8IhDiKIcxtVivFUJWgtsj2jDxNVvNWIo
QbTFaoJ29hQ8JTy3NcME9csYMeILLXRiTlMf4fgSFLNrStQJX59kXTXJ3OhJ8uDuXdmuMoVZ5nwK
UJEBTX9IFHklVMbmz/MLzM33eDUd4AS2Q3oury541ZWiIruA87EuP2kJU5Q9MItKucbSkf4VDCgB
HLBxpG4AyTLN2zfCBKkeaxQ0dd3S3cGK0CoCBZD1mPWj1w7dkqe3v6cibSthA1pNLDKjTuFLipGN
6Uu1QJNqKoR0LrKLDVtG9eg+RjN2EN7J4wfAX5/j6acQHS98InKTBi/b6knRJoo/EADfATE0R+90
+US4As7nrvtyq7vaEVS5j4EIscbTwbePUvqtWE/I2w2nNzb8fadxjWBYQz/U7or98GW5Rwb02Yye
VwjL3EA2ljbmM2+Gm1NYf3E1OlEqL5ewzW/7Wd93rnnGn2oz31HgZ/rYM4VtrPWkTHzKxzxMFUg1
debSrJG8SnOTx4XvaVFL3WbvKJUQucPZvMQfias2yoMMcWdpMT4V0eOCaxwvnGklSrCqhDEtoqgi
NKz4Oe6FGMj+SFQF36jN74zJlgvbU7H41v+91DFOiAEk+aVOs7H+QFOMhHkYiAvcY/bcptZ9qyNW
O0X38wHpYIq1D+gCxd5HZxvILu6StJh0+RpKSoUNGeO+Z/7gBjdsE6QLmDdDemlhKvmuV7btvjvY
Yw98hkABIukoXz9IFY4ZvpKzfe91D/KfCOvSLkorqAQ9/vx5abYjIUZtij7NE7lFJYxTi15hjPjl
KrXCQBq++DV/Q5vGAJNxs8TLxPJVABLju8wIlpJ/H2/9hIxmMLM7qpkGHtU7l7BkV2u2Rh3lSYh+
R784PH7qrpz62hNC/bY92V3TdmCRoqST+IpqHyg5OTaLmGdk9x2idGlBqkup8YLzTeCdQpPsIppp
4/QDItY+z3zO2dkEoj6tj0Ts+5IEdu2Jz9lCpYBWwelnOY/aol2suzWjfsVg1lKYwRtljpFeKmzT
w52pMkvGRXJQ/qucTBZKqLaXiQcxEQLoRg6286ZUdqXcECRvo0QNAbVzxwjQdAQV9tkyu4jmnRNg
e57dkV0D4Q62q8UgSzUyJKi04F6NytyIpR6605hjJLdj38RlNdJHePlHY/H0MgdtKWbA0S0lDJZh
uc3Xj101jvncWYFsNzv2ThdiGAOlzVxvdjSwnru4KnBvGU1ASMSmsdpD0F1yA1FU5VeKR2Kelnvl
upr9jy0oF7XwOsIa5eWXgWoQJmR5Apxzf6Xamj5n45yOpsWcYauslWB3/8xpxoKc/mO+woueGTFl
7klsppYxM1J2pxY6l5PO5dcHzCUxh0iPkY7xeL6W1fdDeTtZD3Z8Yx6hSfZ5Z0sp4q0IGRMbpPfT
mG3geyGckjcyPww6Ai3fuCKhVQlJW3KnCNKVOxqJzwqy9T+7yUB5tzhk/oD3W9tKLwX/joy5O3yB
xENmsi0rg9uHk9/rGy7UMvdU2sz45yGykiCzX9JTAjx9tWIyjhTMfSCZRFPZgo/tY+zH9W+pOR5l
HpFZ1U1XZ48pGAjPqwCrIwKUFvlhngwRQ4qb+1T/+lcXZHZAXoue5T+qhcsh5jt4tFP8Z7/5sny+
JnvcAD1IgZCSbn6M0wbzwLJHAEGS8Ql6yevBDNKPYptXch/QINnW+kPAVq494Nt1/QvRZM9MJyir
tJy7oXqjBOi9jaoBZgDY3eEpspSqimBb97lsZ+TTwRTHhCrT4O3krpYIrcDTjYSX/rHlShINXr6K
1q91YK3KC9j/kpxicZmYTML9BhmHzXhDYXTCakifRtZsIScYv9oVFlif9kfiH8ObX2a02eDvIvqt
EBEbtQMI/8R461U+1/Lo+vw8hrrgexAb7ofdf6IdFrl2/2ho4MMyHG7d6pSOpXKdOi7ECUnouriM
uMxia3ODJ8pd9ShqW2f3j2Fqze9erC0NG2WuBzh7Kn3lwVL6IIVQIMBSU+1kd/ogdnWpsJxui9mE
LHWt7eUzbyweoGZHIMUqSJFQY7hFhszvnXWdslQHs5JI+IH7ZytHCnjzBKgMC8jiMpJvtxhBHLR5
EVypda0LkdVfB3jK87A1cjU7Ruoi+qdUByrJ1yOBH/FxPyfqHo7GyZp9cT+QKKthk6DdpSjKEdSg
ZHyR9US9QLMwK27KBsTSl3Sa8sCwSqTnN7jb7CE4vtjBAZ7qlYTNfRZPrpelyOcYBXOL+NeurdWP
FGOxb673WYLZrK2OcIOwgqAb8xcE0d62XPVc2YsqQASvN1TNfxVPpaqzqiCgLMBJKYQkw5c8TfE7
319YUdnSW+LhRbWzIAfJwHK3bzsMJzDWqb500ciq/5sZ7/4oR1VwgGJBUhq65Vc3H6S38234KecI
jXwscoqac1DpTQ2g6jzMuZfsRDKl3dhP2S0mzMF3OEpY1ugIRbacE1AXeRdzx69UWDIAwj9lA+4Y
hxB9K8doetETnuJX+swMZDXez41uyfniIaFXAwHJTsEGUO4X3scZEc7rspVNyBbvnfn0ZEl+iDBB
ix1Hiv3VmKqi3q+vJLFwCVtmPf7Db0B5FFSDtZGHqZ+J4LfGEEWOpDW+QvNB2cLh+/qj/WwEv1Rg
vZz4AD4GfuJNKIeAP1D3vku50YKYGlYLYv+nTbeIdinKzHh/NXknlWV1AWBMQw525rPJ9sVO+erW
6W+rwc3vANfXh6F7x7z/gFQfXLxJ20AM5stltipJUZfRsxTNn3CupzXf/5D0vSYUZK37Eph1zd2s
0qSnAi33Q1knadnNoQi8KsfsvCu+AKC3VpGGTJBUex8Tz5OysEgigCQeN2VycwWsfm24+TKx7cMk
1j431gCnnyPnPuYCym/rZGxO2SVshd75eSk8kcUUyeevUtb5KHNzSoUoX+6x0H1lwjwTdL52KfAk
N3pOLVmnlRVL9fnlLKRoH8lQPCw8U0Idvp8fldDqcWmWJ4YbjOCTRA7NfLROAGxXY7OV9gqmYmgq
6WFzst2x+kYnlgeHjoHU4zlVGkGRqeSy2C/pNsArzXelXWQpAf0H00YWPQ6MkfYIzUrMDyjYd8Zm
lTEzLXr5Jt6XzwwyMHLVyn4Wyk3QE/aP3QeJaLBT9eqTDdaHeu214U9CtDT70Jz3T7Uf8y6+PQD2
5oSmnJeVdz0IESvGptoKNieWwVjFCBKlrnnfVao9rK96WPCLPorbNiVfq8hqnVPyo63Lfa4aA/0J
mIMaMjFpKfGMLsq9/JSyfHnHRN6qDFCgzaQ6ydfkseJHirkb/JmDzg28PFgKGGTZ7CP50dSAmJF5
Or314Qv19mPhEk1LxtgFpQ4XT76k8cAEylNyhWWfBjlXAxu4j0wwjjC9cGSaDRUSqe1Lb7vgQoQz
CU+BaVXHQguxClsqPUQddWq6eblzP76DImATMzRAFTOWDXwWuJsLYs5Qp0nsiTsy/YBGN9E55ccV
BN3N67hKGxaZooD94MCprZMYqcQa6zrGU5wDQwl2sDigyia21+NzpblbYdfo68uDoVAtIaoIFJJ0
/Ya7nNs3SBv9JWT9n2iTs8PfR0MgHhNX/on2wjwCti3FOHWElFgEk3pWavediIWYUFPXMzbM0CZi
IB2CdyTvJHUpgQDBDzgK0xUJZFxI6LVq7/c9Cl0kJF8RJFn03IuN4AuQXNE0reyr8qCCxLZw4wl2
iX2znltyFF0Da0bOXMMKX0HhVn85FW9qSC0YPtB12OAvZ7ehZUCKJeIpyv6LIoroTffepwIaYH1n
62XTZi1fBdSTPeCZcSJkvXDhlM0l3E8TnVNjIwBVg28TJgzdcdxgWjdtU1REqYx2YmACF2+6M2fX
0W/Xi4FzCzlYeyr1Sq4oYtjimaSDjnODYkIXhPhf8jmiPZmnabYb1rO+qtnDx7M5gvjUGc42abFa
Dy+YaXZmgAV6dIe6bUtGeTd8F3Kg7lumL1qk9kixtul4BIM4nGAsHGXkiH0PoBl2VBjzRlyLiCEh
zl6pjcOYKWsMBw7gTXljutIJWTj1eCjFS0vtXLCaPrDrDE5+N/jPNrfstoQCtYShdf9l+z62YNIC
kmf64axpmIOLUNbTfp0/UuBQk+yV7gwe+IKDW+33SBr+bEILmypfTqB5ECPp8qdeVRlYsRSZ0Ox8
fYlLnerqJuLBzbWIy3S55pGl1wWH1q00TusVOX9Cszyj0LNsiO478TkVnwYp8Ck3IfiT/Q5kCXvz
tCBmur5905K/M8JnKR1OQbNyS63s+p1Xc4yg4E/lj5qP9B2lP2lxwJ09puGBEgXWwt3eNKTdnzdk
YDciEMGmZryy1iDfajrsTfk7mrovnAKnSLasDPB1ZDILkJBb41piBC+cY7Etw06hDnzh4jXWbkS3
H117xJq1P9GHDOfldHtqPbIHxzRTUnBhei6e07SFi1OW+4eufJHyaDPxiL/8Tq6lcQuZVRaqHk/n
pvReFaG8hVeaxDtF+TZrKWKaOxXvask9R1+Wbf/2K9Q3Sh8I9PNM6ShtKSt2eztU511smjHQ1JSk
3JiCedWDT/kHnsa4jYKOl/6FiF+94nGPMfQ9ZUcM7c2amBbLjYSDfYOl2nBMESDSfePtkIuCtWNR
pToh58MsQoAXAyrgn11ibKo6qMykAs+Gx6Oo8bjDjSAHEyEnV7hzylTbpaQu3pz/qz29Y14ZCkRK
txMyPwSVyxZyZyutYqjUUdL/iWLjwHyiBVGLUsJpmIjAf0hbwGeQchUMNeDh1LLpBCX5Mv92wt9c
osFLmYHf0kMFWkKovUDIAfc4Jn/TDVd1emVrJ42smc6/diQEazo7QwJzygxv01OA2J8AESBBQvo+
IecHKsowFLreqkgIdVWkHEu+c73KWG1ZROL8db7p0+uTwooFptzmXgThEAIuCraEqtCLrED9dmgk
TiinDnK4ewq4eW666lEDNPkAfru6um5aLOgRJJHQoCSNsaAck3Oh3c+a23Yflh80ho0gO6cRfSm7
5Z5CTuWmehgGBSU2jOFSiA3o64KlEoD4Y527vFzsj4QyMf71BIrh8cW8iw8iRSbKvfZtlqAa50YH
u0NOlL+if05w7UbrpCNJUaHUGbOUyG8/GGU1k2ZeNZ5+stARrdrOa0eNxNUvMC1GyMGIBpAzTHAy
S9lC2j17t9YtJK2W+Nj2a0t4YBXiYUaLq2MjOPnL8FmVF0yVTHFjypyVHPPSCRpJphrKwzfM//55
WXUVScZQmYfxJCRL6IV2NvGHaoMoNd6RpqTITDWdKyi73Uih9xI082Zbrt2FAwC90iAp9tpoVUZQ
BTvzG2s3vIZvRRztXYaJHbVN2qdV+QxrfHBVscrO8rYH6msuc9zkNSKWKSKpTPwDjkBr8wmCtHmD
7M44gaM7Bt0TFD5A8zkdEAd5sTQ/xSl5VqjfNqaUcm3TCbpD6aiYawV0n+PJ4lf5wb7C1AgyWKLL
odMFljJvbyqashKxaOyr0dleuOx9Iqf1HbEMouTu9gbAJ2fZbhQtZLukiGyIbWLR5rJA7RzyC76y
l0AAIfN+Uhe5HOhCmZyICy+Ns1ETfb2CRMacfSCaW21PHKXCuo4cd2enbnLBQRkteqc1nRn1VFuu
AIWmMnr9SrLu0DPKmSgGlMnfhtrnjN9dyKWDBWE/kkjaMkid61685ICF48QGL0Y/O1kzlYUfIIOT
o5oOYiZOxa0WzsBVuLujUs5IegRBg7TGh6m3vi9cbp34+z/OC02cARJ3wqx+4mnwuoHQvu98V9lv
ZmC+zarO9T0IDS1z7hBLsQq3gs8W7N4154jiOEw/dEYFawVDfh02ZJZbJHnJ6B6JsJUhmA7lKP8G
5eLkOnnTEQP93fPj8shyPeugQEoqpW75g749yE7NKJCjmLTvjkS8VNtfMbb+W66RmQIXgXhxsCbQ
7oUS8wqSv7zne9dbSP85jrX0/3smi/a/U6/6DWiDdgeh6mHuZWZyet3Ty4dZnC4MdGGR/5mGlUKk
alqETuNKd7226ZJATXUKgid373HZyKfZd8vOPP04F3mCrGvu8SDc9Wh2X0KLiHZjoRkDiuyTCmb9
kroyUPOgXwhbyHTh630DqQO7VaLrYgvzXx5v8rycvavjoX6sSCychnA/P9Ej9gSfO5pN+jMBckoK
8nNZta0JthjLgcW6wBtIfLMKa+3CYBgDmNDOmRvVXCDpT7TSMz4kB185eDtNhTr8omFSXuL3w9Sr
g/S5B8P+0Cv+QKqc+kRyZnOIBIdxdlLrm3O6wSmGrNtLGYKkgJPaHHXgF5OmSNRx2gtlYAh6YC97
VO0TwwsbFLURLo1OAgLfkqNmocLVjLjg94PU2hlCGc0MdEwyjSzdp0o/awpJxbPUnayKSKdQ64N5
lI7rSrOscy2Lc0ihTI2+Cw07FQ+6yCTL85PGf/8NW+HMofRYPMUhOhcDitjDI7RdHAvSbY8qD/Ru
qijfOSa0GaoRQMGe4qSVqvbZfrT9ofEXTY2NiQvzMk3cMwHqUPTS2cCFDwc5FVQVHwfBjBMxO8lV
jFV3j+UW5cri+jlsZbP0psIFENvtQe45z63/reZMjW3MosKXh9svQ59V1YxoV/NmafN1gQ4dZmGA
M21UwyLoCTExCjUXZrvBzyumn/UdPbpegJ4gAzZSctWP2Yj/N9/oeRmvHcYDUQUK0+akACmMj51T
5q7jAWAaxQK0ioJmF9ouqaWmsN/Y6wOe6CILn1DYdy7ADr0naXpTY8BNRZfX1GcGKHpaEnEXWNJT
nyxAzp9WyHl5y3jT4f9MRQV7280h/WwFaqVkNaGniueFXJtIqwXpqbVy1Kxi2iKANgfxNHbCjEqs
6BCizPUSM6xYH2dQM6WnxDGh6zrxBRSFZfpsCSPl7yOe3NbN/aPuXHrGFPyJHHsgKfwpPFcBVvXu
GyaWz262nmeZipeS1JyLM8h/iqoe5/7+vIK9+luK0d6ikyKa0+Mn1kDKvtc1Xl9T4C/SUShnR5fK
oqJV+Qdg/2MpJ0gkAh1UVzjieIejud14Q8+iw9DV7tHMVT/UvDo4w0V4wxLzNd6jszh55acZguFN
3D/8G7RHgKdT9C5lTPo0iDqY9jlG8+ewib0r6q6Szv0FnO5D4Lp8xHYwFVu7qWQftuS/kvxIROec
gcyxURTte4TAp5DrKptu8N0FuDnWJhHT01B0xa1yRPQ2ILj6C1m7VHaMkkjyey5uTBoWgcqMIIZn
bgBZ9ATRNu7Tx1XTyjT2L7KJtlHYrVhps7LrXFehqJP6iH9Bjy3JBj6ewrttJ3bgmiM/Cwb2An20
Aidab0f/TR0iS6NDTFiJGX2Gq5gag3ddpHNccyHXyOKF1C+LrmU6Qf8Tc4aKs23DM3qD+089DdKT
nAkbd2tJSPSQqlozVo91ym2M0Rp+Obw9WNglUd80l3zEmOyFWjZhijtQKNu6Bpzw1WJYQIOkn3/l
L7nqxCxX5WVmGPPq/7+1SjXteKs/NQ2ahvBLyuCnVmbCV0pjZq+nt0g8or9HIqRvIfuRgMVfdWj1
j99C4si5oLPH7QG8hOAoqb8IGuGxcaFidwGV1gBbC281sdq/KPo8o8G3Lz5PJ2XWb63z9K7XsYP2
Udo3rkQIcBR4EVcTbRx5ojy1iMsQBYo2D9MwAJDm7syWH0kPTLwfafkEmiloZ5fNXwJhAU1gcBWF
QzHcJiYwgg4UbzX5Lz71CCEMR6fIoLGV73nyzXUchhC3jfAm/gOTKHR/QA/y2edh/gpKpWLxCeAj
FF+rEVUTIPLel5DV4oRuulZkfCdiJbPpbw5m1sH1qGc+DXf+9QiHOIULwZItGlnJw9A/WUEM6UFe
PItYUppwzinBKTYw+MQ4QWp3MipvAC2YQM2IOBuC3ehg3R/KROyY/1J2rSVfhfRiOSZcFUxoB5Vn
lQFse0Wki0uwzXrw6qog3fcZAAZAl4lVYivdN5J5/busbxV+ULKu9oo9dUWl2MtdtLtL3dOSCD2q
PwVfLLHl1ztmsnlZ98MH/wGdodYIzvzH7DXn65eW+hzgw2WznUf47uj+EiL41oZ/eJ1LxINSJFdX
tQoJZfBR6IqD7sVLu7ouaB3QMHTkGC/b7s6PBJ18HuBJj/dn+p4h/z+2nc6EZRXhk1BP6Gfg1Fwg
5hTGr/2/d8iT4IfocHzpMAXNsfiVlC8ELYNhSIqgjeWuYKbdMhvdxf9zqexwCuRog6x/XrzqRcPV
n4j9bJrBtqAyGa0Ix1lGFXZXl/IMBwxifgSny6W54AOP1fZ0qDTGfezJcIU4eV3j+Q8F1sTFEQCC
fnz3DimW+L4dBQwBqR+yhCN2Qz0Ed61zjG31I4m/rJ5MHMMdUWBLobowbLkS6EdxqXvZwUO7iZi5
zitM36hHCUvigrV4Y3iIf0T3sObgKnIb1dGTA4Yd3LuRYJcxzlezWCrN4L5hJFWkocVvcNa1A5m6
3WaNIPy2g85Xsce+OH5F02hOg61PmjBF8a/CQSCUxezJ8b1LGOg2sO2/sGioATozdfrEgr8RtRux
IwPJaxz2xxl46NOwnh4NwKIpUmgmHDdzfLEPK+6oTmpIPCh75SnwAreX2vQ0VBkiCDLleiuei5zi
NI8WyTRJpVgg1mguAWLOuwB4ilKVNj/SV7L+N4Ql6qDD0Ja23C5b9URCAVeeW7KSiuKKg0wzlw2T
JIz1MzZ7vLkHBc5YsMRxndIRDYbvQdi0IPecZ5mDzWRoL/pMpWT7PuRDZS9w4+afHd4fxAsxn3jE
5CKcExpJbjjD6rVAPYKB1vu7dSytBdoKNQHsT1+g9FbOrRHJajviv4uIpE6pYppjt0O0eyUO5oF8
mxi526ZJowDReJH+mijw6tm4eMceoQhr2J63heP+HsFx0g9GQagDzdwmiDyjEVfx4DwHmio4RBSq
tE3wFszQxleZm+Ih5H2JU5jcu8WMaiSF6tWOjBGhQWcpy0f5h1S96zTQbzw89DmacayR3Dgpy98Y
GG4aaphTMt9kqUoeM0YTKXxEtOgr/LtPF5XGmekiH0CF+UDCYfc0SoVEcQTin0MyPPw1wrMmqVAT
YtL3HJwRW4t496E7vQLB9ho3ukj179PoZP0uuRhQv7VuKm1LCE+cXS6w0s0ChnmjURQ51kkGw63+
aXOuBxxjD665R+XMYaXnNa+ttMbk8zr3+IFrKgU7dyjd0AN2ew7PDzATp/Y0dWwJljPi/P78vYyq
MCFMlOOk0cv/QW2JdytIX75lkzSeJEzy3HBiqA+Hcn1sgRsF14XXrNSnH+IZZvkxj/qmmeQvjEcV
9x8kv8UQantw2UKxSj9XBB06sKdO7e6F12SNimD6bCzKmtdYzZCi6AzoETOv52eqL1KXslDaIY6W
rScMprgjQI8LBlGCaVVtcfq31bc89d77Z5nO64ZLuFqgdabnvalY0V/ZZ0HX708u85NrzbSNsOOx
/oKleNt3AA0kmQTZbc7mo67MauxqjU9U7KmBlBFj+ycjwV5QJ1EMMhwEyCrtXI8jUliEgzv1uQ4p
5qzIqMFIQY8/aA8NM4d18R62EciP63GyK4Ll6wOHvcObuogBXaPWp4w6yBxA0wgJ6ElOpUcyy3FL
97oqKymU6jMX6QgAUM8uL1B4P0/H6DvHGwNCW7gOEoJ3HESt/VK6DKuE3ltUbOs2Md2sNn8nm4l5
s58rnbvAd2LGSWLG6clf6fswfc1WuUMRIDfYeCGaQ4KlvS8k6NRJpnXubZuMLkA2lkGTE3vCN9So
fer8ST6VUtxiaeOuPtupLgzJk3NQzUKM8BtNDUGiSIzLrpr266CdH8vs+pVYMPaGF1C0qZ53N0Wi
oc1v/9Aka4z3jVb0kI6vdaFZ38FPY9c6/NXGiCvDwOjI36094CrIgc7M4O7iZkKz3kwYw6W9S3ux
nDvrcW39l/UEpCCFMTP1f1RcQv2NlMAgRnt9k4u6DqZxadW5iHgfipsnLt8FgMR+e+7JHCPB5Jam
2eKkjFOmtGw78H0aV+nb/M9Y82ArkWyf44dX3Jg1NJ2WUeHTs6TWfdPk5yngAYlEXmK3O74ampvH
b5dllkI5DIHW4vojC0eIzpf71fRjxsLHY2BPWYcQiJnKD1dK7bPGB9BMgefqBxfz79cb4bYA0x1K
P/7BB6+Pz1yPrNCvvK18SZo32U+yB+BuE1g0utVikyJVDbInf/4bRrxg9LsEu1qkRsftG0nI/j98
CRwwC5c3JXV6Wm5MxyoHiSOoptYfYKEIdWepa09asm/NCMWqd7B3s/wPwPrNQKGdhoSUZn8woLNc
qWDcaAveWcqy/xFLmuoqbExJXgzvvVZbwTxXjTnhttFjCFxJ9zR+vtedn/1z9iPnhrqwhn5Kp8lA
r0/yngyxjx9Uoxk0ENZ5nobHsXveSYvI9Fh3Ml/3540zn1ebyH2Ub4uoQ+kPTnKbFnxQUkCRw+rX
n0eOfaq3SEpNlcJ286S2stJa5B1T9opDkacEVqyf/bQ+eO4RXxm3CGjPLSG8bcpianHoGd39mZSR
Bk6Y4QcnQG2/fhnNQ7jb1L9NOsYOxVdkiQ0S40X8sAbsIcZy+WoEvhnKPF25isirvtGwEVUUJfNc
G6johhY6MHYsELC/yoVAjvjH9I59RCCO1JUda5l6Vcsx3FwWW/Zp82pPXlyHnWeiD3HbPoUW6pMZ
eV81qideG69/nJEioDZExWb4aKZujZYPEEmy8y8DxYw7P08Y6pxjrsYpeVV2NbqlU/t8AUttu9Fw
i18O3qpvw+37YjKZYSQBUN4SOIfcWZvUefqHlWZwXkAOkuwwup6NFll5ff5+Vzr9bNOdcSoeE4BA
At3rM01KFwhoaaeLn3rssILuLZHuiwi/PvT06boCsh9yKWNLtqebtzBZKiBhmeDT4PcULpfM0c4d
V3yOMzgyDFk3AlJCCnXdXNa5BXdVJcXf/8+Sd0E7N9clIYlS6jZx7SjpOr1g6fSaCxzpqCmOPfqr
4iwwqItSuZuCs/9w2ddSfHKUMZK1DjtLRMM2M74yZIfRDD0mP9DdtUR/Pop279qGoVV8yYflP7kn
ENKl8s09s4nUpseEOCBsG0vd8pez6AbEGy5gtdMjkoJE3kTcycrwDknhXb0vGjp/GmQV64VufhkO
5VjRW21tGOSODw/qqTdFvbgWA6tgULpI+obvXzRqmUnaDn9W1VB4gXHgDvwXN3WuMav67lTEi68/
Y6tR9cA62iK4PRgWRoqKT1kfVkfRoaE8J8M39XSNWBI+0MG+RzZpSXevqh1OghseJZPvxPXiEuq/
gbXlffQs0Z0M6XsIaAJa0WGob3TzkcwDvCnj78XYBnWM6ZeZ87w92LAgOgOjtpwrMqeG3vNlE/aE
I90+F4vOoaqR4QXnY2OsBywq3pB7T4looGuMHzRJ17iyK+BJUQ7aZ8Yd9baGZIs+QWSxOntMvK/9
TxNX+4ukFpVzHtYK7BOKHnLcjV093KpwzBY+gqvkYiBq/cZTifKN9HuC0RX/eE6duQQQnf6oFXsz
a+0DeZRouI5ON8n0V3Fuk0pRbCqb/1m6kQCQejhT15YlyeJkfW3252hJ/Sj2BIlpend8uxv2Z/7q
OiKWGWNxQ1rO1PFL/ZFguXYHruXFwztXROdsUMAp0NuvJWHlhII3QT55fHeP6qMz15fIWR5b2TTI
4knrGb8kIheLNVRGHQ3d9mFMpPUASQB/Ukod12yzWw9fo5BYu4DomTxri591pCWh01eAaxHDOTPW
hcvDV0bxwzm52kVL3cP7XkvBfMhYXCc/049KwhKrJ4BNsBKvSxWmrsPuk77s+mGlnB6JyG7DGQ7k
I3gLDxJLYbzbjRMCIJZ3AleZuFO7SY+FNknaBZ4jLjkHxIBU6MOO2PAPngrPoP5kwps/Vbe2Ibo3
HN7Gjssrl9/b+8ZS2YU8v1t7Ajm6j1XJL4ZE56sfrDG/ccFPEz2wd5jVAwhkNCHkbmTGejNJTb1U
4965rqNGd0iLhq8ZD2z/n7V8hOwWBMHGiZIVXBUszQ9XDCi4ohmUuDIjPfMqeHO2mdJt1TCz9xY9
ByCOBHepoldvb4F+ME+Vb4/oJBjCp2jiDRwNG0cy1X0XaVUjQiy9vQKjiPv7iBYwAeQUoC4oHfzk
BtAp5/aPyq4WMIWH+zh3DE/nWN/uOeyIf061U+03TYVD9yBCg2ynJjBnAextgmwfd11Jyv7W3bkQ
YJyvE0leO8PY1q6KJIeWjgnIpDgw3+PiIKrQYReCYH+KKk4x3vB6k0aHq9cHrAF+UXvEU+FcWbgR
pFlje2hi0yvtzXTiyHdCKX0nJT+1eR3uBlTGhuws5bFuU8ERT2KTX5bzhkcUpRWqNqn2Q3R22WsU
0Sg1Ra9O9et/ntVFHGdYg8GQ9oOG9AHQ6NV5cvXmCgcWHRnWRPs3o4mQnbly/KLtt/UtACeV1Rur
T14V4i9tDmdcLAM5smfGrez597+fxX6mvUw/Z5bOH8bNG3VM4rPXTLxzMJELl9kuAQ92nikh54G+
8oDicNiMJxeh51wqU+y6/NKUQ7tEnB8Ce3CxmatI2djtSxcuCLFqmCr4Vxup7szySKl7FnCWgogj
d8kSkQHzWS+U4Gmr65YwVf6wYbvV6S2WHNjSJj6I5fO+qH+9qu0GJEjq2QUg+nrfiWwcZo3rwV9Q
iIZ1O1qfyr797dBL6kH1Aq6nxxOJojljtWft/VGV297uzJpksHPMESXXltzbp0Cr3THn6phfevv/
fCuSclfx9f6tCfWe7Nn96iP7V8SVu5XT4aUgfOpgXkemA/0Gc8ioaShl6MQC0BzV6to5Oo+Z/ayY
uKi1O+vTrnkMPY+d3F6bxaVvfrQnaOF//CDZXj7lHaODgVnZC8bUEJkjOVpNQVwiL9M3Fpgwn+K1
loEFPznAGoeUQwiuGLwsnPdYfaT4ksJwBUi4eJL2CFk2UzxF//Cei6JmHFEtpjmct3qasDwqo5IT
U5jcd0R1i6IjCzhXWhTXe8sCJ5aGcC59lFXPs2qfSI6ZC5jwNOoz8wik5hUWoUxkrkS8Zm2rCnqj
spgCsSce3HmQzNY+5ad6/K10xMTq9/W7qN/n9jOVHiDGbE/4V91l83Gk3Gt90/ewI79iZgQqemW9
LEX4uuFBFFJlc63wQ1uAEYTXOdW7FIFfTdCGUQnPAnzXWSbdSNAwQSdgL8mse/AFZ3Wbfqt+8NIG
RuP62ZKhlbfkpe7PgaKcyh99yODkovKM5/wIERwzgiR6PvcfSQHlJ0WerVGk0D2xhO8tS5oaAHqG
ifv4i9PSUiCcZQBH010qACCV5LzPpQhoiJXqQUGMn3hZYITxSVArlWfIapgjEfYoLYDWFd9sqSIt
lAKVGcQP6PehaEARQpprOR5ujb1c5Ow/X5LAQeUh1lPtW2pE03umgrYK2Tg00XZogtjZPqhD8RiE
/q5YbhubsMAi2cshFFFvvTsVLDfpTPDScbR2YQyasSG9RLqBkavqezSBWpCeKrpc8vF5S57/7zmZ
kUsfHdLkPhqT4T8VVAAocvYJJvZMZNTGtCnB2mx7xTSA2iqO0qhZ5Tr57Xgw+4cnOPfWl0MpmZAy
CqStx/VEezWi0JMwM68CgD8NpzR8z1Av+6z1BWUqwDv/d9sbnVVclsNhI8c5TUCOx9rwheS6rmTV
QZ8ZMt4RLBLrKd+Tin0e7lkDrtN+YKBbPzyR6MoIbGTS0u0dWVF13pFvjkHC6hTlBhai7Dc9Y6Rj
e1QPWtWMcBg9xZoS3tcS6I6GKh1YsDrAIGlQKHvC1gBHbyydR14IR78CW19QTT7ajNvTovhojMTd
iA1c2/Crs5Cl40cKxsLTmojVwIFLicISWebcnggN/iG26hlknwil4bNkZVNrYGEyF1d1brhxNZIy
M90Cptqp5jsuNIb5LrpG/6XNuY9Mly68/MW1+5hGUokkeZWdHSG3fEsLdgvOtey8fX5Nt1vPxrlG
RhdwSnWXvFpBW1Dsolyfc3iDiu7aexMM/Jr5to4CWMDdKZhENTlzpeQVj4OcOG9Rh43IQrlW5PWq
Z4nDrLvoiCtz2G2J1RKENI9+D3ed0NPB6aWZ1FzJlV/jhwGZcmB++L4tGa4/eGTUwV6LYv/JEJoM
H8FoLvtt5zChHKgaMRhg2ONaWgtOhX/imPkILkzZXZDYfksfAYPSkrq0lg2BddI0xGkzQwXl6DI2
5FQL1rPLe1toy6kJ+w5+jZdH2eg0OK/gqtiFMJ5A3zqPXCkDXvI4uuKixcxscH0zyv5j5fKEwxLh
Cjjz0AcpxrOxQGtb5azRWF4p1OMzf2H8wO+MqGfGS2CFCTjBpO50E+nv8STZzrihSBn1r3DWImLP
ZqTjVXGqkTTPSsto5WMyHjMHUeVLzvxfUaYhmYfQYoTuGlSUZyjKcx2+o1fHzA75WI8HKYKheSw+
ev9DL3IVYcuWixM5sNzcghnqqfzPDwSvkj84ur3t567KhqgCQfv8vMLzr4oLByiFyE7j3bQTVcPL
dmkNDQypPKzLJZLICExH1kDOq9dPpLkXoC9bGlAnhVJ5bPu/rdbxKbZVTOER0douid9nYkeZi6nZ
UoxrqRxMxhVZTYM3D1D8q0Qjw7/r8kdmnqwWiVwEAfbckct562llpRGLVNTUbo/JLDJ1TA7jLpfA
faD5snBgzyke9hl6Rwt/0swzhgWSJfIiG75wbtcFDtyrF1hjSWXw9XkKTQsInWJjPT3LdlIq1UOZ
GLB0hpkEcLzjO02f/LQ95xXxnhH5hsQ/GU0QcX+LbOkU2IzJTm4IplCv+w6G4WGu3tHj2DZ6QA6z
pAzPX+bMSW/45sjC96PrLn//OJixwnk8RTElYgvfezXr3PW9O0ADb4Ghbmiaw4xSREs++tT5G/8A
GnUyh2f+NfJYOnZbqIKHF9h0WPF/ebDewVkg+JoBG8NsWLBRY50r2cajA9mfRc1+5iMXovOoeNZ/
97YOV/vqOB9JsPyP20woV1p9La1dZf9sSheufCxyaf93GTUEbFqBqw0711dIpiZHeMsl4cZV55t9
m4JriYiZhBq0qw3kDiXy+C2RTjY79Tnhnu5DQZzybDse1hDKCrIPKCR3XF71ZUI/+CmBy+pdR+N4
xPjSW0XTmOREHLX/9esCmyXpJoxchNqiCV267vD/6a9yP4Xygr0l9mnyQfvW8lSzs4BGMJdKQp0h
01jSyck5SUiEvE3Wiz9JeM5U7Cer8OGxtbh/DaiTFs2Nd6EcglVmVnc0xIktwAb7E7xSSKt06cPU
Y9sDp1my69JM05CS795ErbFlzsgrMq8IAt4l2osiD8YJIKLI02E3qxT8jPz2RsnocdV1t+IFF1fx
yvHgoiDNr5SV9hnnsnEh3x0XSQ3PX9cKwwd5Cat/4IC1Bf45Bqhj76SgKwDHp4vHMY5aLpk10Gm3
iTZX+V/j7slK3op6wYfWtxgoF2+7YcM8RJEOzyEY3OM0TVASN6Q2JUmH2n+RheYJym5QrEi1h4Lw
R5niJsjQ2rzh8pRTDR9gP5SH5noWKRYcRbpgubdpE2dxBq72mRlFPLoJBIR7n+9cwF50IYJbEJBd
zTslXdj5dj0okIcv1Y85JYe6Ji5ZP5SPueoDkS9CUCBSVHsBSSciEk0MLIKfY5uOLo7388jmlZ6i
fePb5A3MbT92OoEeTY3zO0hvp1wi/bVCTytrvYw1U/zAUdYsJRIm6z9I8YfeAj1b1ljfOyvEDbWj
DIG7cxUZzPHBshHCfXZW0+Sba2tRvJ3rpAEXCoUSSAqdq8TyqvTDCwW/9E4yt0FTuvrMzWNZzI3Z
cJX5ViXaMcGgHA9T64ayYe5VfjRwnPO6HMue9hEjrWxs9w+ppAUmyGQFYSO+35D6Sx/Vne0MG9w0
7M3X/xi2dJ4OPC4L8fjfid0ByKZL+6gCSOqYPb+Z3jl+Y6TOIq+pLyTUOQVcKShJdvd8NqaQUvai
h4HtkDdAQt59nNGOFJmTeWRpMNVjZMx1/20UBpkEHwHS1tO99qoARvyokuqwC5XsVvY8UrNIo24X
ULUseNqtBh+eu9nG5Q6xjF61VcRhAp13/9JeyQMI+lh+VD0k/+qW269XBKTQaXzRcrf6TJAkXBAJ
dA/BIOKsOrvONZBV5AXr8uu/5MakhQMjWi6Kpt22z/nNmRWhsKAlQhaZd9axVdSP3rgAec0yWuJ3
aaonBoCZwtsSDw7kgIgjL526axq1oDDH+3fm8ZASg4ndZ5HJKryoj3s2OTnTw1MbW3DakOl+zI/a
UyfO3CfagHhxl/gemkyDsCAfz2fgpzNhpLJJ7DLi+qG/ibarLTm7SQEFNensP43QpToAZsTqLQt+
S6oz4R4lPpLWdT/A5PeVmyFsiQY/1C9RpaMQFoPuVtNpRooVpbF14fPL2r4m2BR44FA+tvUJaFyf
EtXKx/24Dw5iigh60nIA9wN1ZC9vDz4su1YMUbKTOzbFM3C1uap0llCvLKu4lDbjC3+62gMGX0+Z
zytx4GIn9kjtlkJ0N8QW5q5IVSJW6I/hHbkt5Zj0Pd2+m8g6FF40zHQjVN0k28PEumFfE7Q6l2Mi
MtYvE3CHKvZNOzy/+UP8FiUKjBlEp4/JNxftqNAOnCcuY3sCoQ4DRDwQpsX6CK8SQL6rCqlHo5i1
eOdX74fZzcRRVWqKnKqpj+TNlp/eiIE1d/jcTb7BE2xvOZQne0rGsd4Ly/iZofVjI+NbGsJhRpf+
ilvelHTI9eKZkem4qiycgnAvp+FpdlGNbpZo8JPxkbYPUnvac05+u1godvMsj9Esk+fwzUmlgb4f
DTLtyO5fHGIKv5S0TrFn0LDsEA+Ylj0XS9H4FhoJiBiGak92BKlYboM23uInb8xXVc+Bu6fGDO7Z
mMTfCtS6w1sdCpXIS1a5BW+UPk0MmaPgHpvCAiriurzpPshuffIOPT/glyKrM1Kqii0Gid2vHjXd
oYl3oBNbRjryioMFBTINutuXDkXworHqWC6WgzXq8RkJqwyST7Y3xr7zZRd2YCPojS1nRLsPEqxc
a30mVVYHfNobbny1prRKLLUc+QW+sFTqXjpDpdqLbKrjSg25CHFcRj+h0DN3nLaj/JpN+3VbWuc4
vAiVQgA9CrjLDI92eNAIyJ8CrYn5u33gQJcEExY/ekmIls6EOnwbX9ppmD61VnJ3ybE1nqtlkkmv
zymf86WbqlZvL0sGsL53WwPk/zbt3TyK9V4iJ5vWVY/LifzITcFZVxMqN462wu5pTRQn/Zhzj6T2
XsGD8jLY4R3wMd/Zzecs7iIplcL3WYz3GKKx/ms6xxebCzdkQi8izox974dEYj8/g97R4SmUpQzA
ndavI/XQd6om/UvLKPBKWwdyEyyj7dSjGdHqGbfITr1C3zLGG2zGqWvnFNt9/Fz1BNzu51LZf92j
0bDvh808AbIL7ccykFeT3ar3PEaFh5MbLzhBLI7yr3Q2QqglzKQb5mWox1JB9dDPJ2AfQG5riSdX
Ui4bRvMZ4DETLDry3qvr/o6rXWR+XVjyssuWllcPAosMlQOdSKTZYA/LVXnEzag0aDTM+UE0U4Fw
Prr93oi3Ya54LPE4zPhCgt1Kj7T5mcjDdwqnwAU82PgW2Isli7uwqKdM836uY6+/Z4a2tMVKDk2C
1fjcV2KGpKBCQE9IX277i9khCJlvMRB6r47F1Ezi+6jCKoNh0JTjk4cUs7FSukBiD/EiveBAkGAV
ROQTsUnrPOpBVBhN4IDAHuoqfN3h/QCv2yINuxLGnqjUeS1QsL2pn0Wh0QUtfDbp1ejKeMRT+Syl
cZ2FolwViZxRRKNpZ24/5Edc0EK30ZiEqW/RUKFaDNQgRmPzIYX3uv59lv/qxr7sfIXer3Di5930
T4DqgzdVFJ30GKe1HTnfW+81yLAHPMEKH9IL2b8tLmSzx2G5W4uwBLser6gTiOIEyKfLSSIbfQ3Y
7xzIbvlYMNXrqf/zPIV08zbKVlfbA/nzCqgNaP737u64kNSqqxpcumNg7IeXX3Spkqn2VOFhBtiR
NIgv3Qcf/6AfJoleNxItesxrPGWdmIpkB5GHeoYujJphIPbmk2vFpHZx1LdwN7sjg+555CAgdG0o
EJxqWI4qvhxWEhDdymeU38jTyxPlpBHRJjCC/swTzvlqrDzP9hZTMCAIRu8bSTK5LYyWgYMNrhfO
Fkd83Hy/WsoHsL2z/Slbu4bUJ6dbn/0kgjwv4Wc1aCmmjzjxObjnxgd+CZH24RQ8xssPc5y1PdNi
h5ihpwmR4iQM2fWhbTymcxJTZZUFN2n9VK9LsFZqs+oZaytpG573EUVAqikgIDAtlCN3rEHjFFOk
WcFSaJ+af8ZEIJkdpru8yRz/PuKLJeJKONhMvI/OOQ/b+Wx+RaR3crNg4ng7nZBLWRasTsIuZ7Q8
JAV56eAwkRI1k6Gi3r8KYHozSp6dgiHa98SNokGqOthscfu7mDagFsi1LfAm4aRxzCT0VthwwZ8g
Ymo/OpMjxvS9E+edcfoYK7Z4Xpe50nMrlKpzhQcMYzB33zNLMob7hvRUKTHHoB6ngIB7oZtAF7zG
KJrmnhMGiKjp0WDaWEh72X3xvkXIXepV7nR7m95mjNIBGlgs7E7QHx6lHNY5rMFyuSNMKXFDF5G2
xqZWsityYPqV6uilnXqaErotD99mnRv0vV9mnnDjecAPS82TdkkWi7zejk513GtE4xopEKB3tDqB
1m8xzoMmePdf9hRvjJ5eMEjJw7pP2g0yaER/Qy+okGNm5orge9jPxnp6IVZupJYNAY+HlEPUTi2S
tsNiMWCrk2HdAQndKMKiniCA++DJGaf8H715aL2XVgJ+WErtFsynehDAMobFQ101XljYaiGy5mql
dV74hUraRt5BiKx2s/KScdmA3HErFJ4yziKBUKldapbunaizMA8sxxQXiqoTvWN6bIyVv762HD1C
fTT8FurichjT64cusI2mtfm1lF/i3Nh+BsYCzIFpneGssRnVZ4mjBnoURzNM3121TDUoe+UFL+Ih
7XPGHrZrklHsYgHB+XOaqDZ22Zv1Y0UJj4xLljLkCLB0Mpk8TO6wano3zVEf8METpbUx4hI7dfsr
wHODDzE+9ppWIAxUbppKGt2ejywZuKD1qDv9fzLRgtJ7DfYJchY4DzBsQ4EdK28ACDZD23D4on4E
nqfIDEHb+QlludMuRya3HScGSrTXkY3xkjkZAQxKEXosK7zm2+15nC9hqRDE+W070BVTHSaZl6YH
PylGN/DNoaygcnS+1XCWaliWU7POS9gC1qcD67QvEZ121IwIo466d7auflPZi1os8kp2h/+vfI0G
gS8uxN2Un1z13LW/dJnPi6sgf8Wk8Qm3eFjN3BMux1NRMHVxB5wXQcu79D7A79tnhVzQLMVwdVRc
4MBAsrajPKdpncC9w5VgmlV60OeE75fQJ76s/H4oJlhpY+KoVIGLkNxCdPloOJryno0MTUv/OjHf
Xm4EH9KUtg9MSSwCHY/xHKPoDcujY2nHRS2arjqSaoqd5eCqREJ+TpN8AR8UNPE40Im/DkA47eAj
OR9Hh2UP36FS1/D/XdqwbmZ8CsPbBBmvWYOCbXORiR4q4ZBGVdwBKHfEmk31dmdfrWvxDq+UdJAP
cihYgiy9NraWX8gKwy7lL9HVoyJ/3Mv7S4W1mUd/ABghiLvzQ5qo1nbJa4HJspDEJh/nWSWj9ZT2
YeS4IF57hA7Ei4JpjprBaeu/YkFzXS2BQ6UUJWCK5ZhDVA1qaCCgQQ2qwNXE5YxGQVw4bgD1bsNR
GyKmHJP40sRcX9hdHb2FUtfF5sXd1CoZk1Zzj23xC6qW/n9YpZXivZXngK7xKY5Mb9A4cr9qMY5j
VrjxZ7j+smT+OAgyaVzzUat5MAqP7l5/r0Wk0d3OCczMy7MyK294iN5ufCDs4Qm6qaNI56pLHIuv
NUDpAH2deXXl5R9j0ZnU1M03Ml7OOU1l+82O36M+M74Q1ogTnl6RnCnvUC/rzuxsohmCOLxbNFmi
+N0y1pbmcSF/7cZ9FYiejb7UYgGcA3LWtktnvomckQ8a/biQt2sk0qgdtIOa2FjYy7lwx9zWYN6+
5hj/T/OevAWpeqmHnEqZG97QAnUd0YVy53nR0HLyDm9VR/1/u9ihrEXLDATBfbbVWXq6Z0tgoYAj
vlTdbhMc4U+BCW7/0Wo1zVvE4h8Aa1Dz4pqaXB2oMz0OQYXjB6CyrJsuecmP2f97GK08SUYdfqnT
UUeCpxkDfuyYv7B/OThqmV2G2bZnOLYP59SAPSvbNGd6o1EKnsfxSysgW0u6l0f2H/3oGlmszPcN
UKD5VHbfRXZcel19AYVu7GZBqsIrMm6lm0AP0+pKNJJPqTXiG3QvynUqeyA38NYhi4ysAz47VTdN
0Mgz2RwEx5VI6Yv+kC9B3s76vHdTPEnKRwnnHyrEferhbD5O4iaVpcIGx+kCA4RaOphE2J9WsMag
DngmRGSXUE+NFm4184wiLvbdPxOhIdIkZePJu8QOQg6ZmG0qF7xLGheE9mAaOMSGYT7XIPeHGlSG
bxhQKYJceSCeKvWasTRl++f93EScWmf2eTvIQ13sNUj54UDC/Zh9B5cp76VE2KH717gSc+gIzX4t
2ItB8eMWvUGrebZFRrEFE4JebWrxE7UUo2Za9PUBGx1hvqLtnVFZWXDnAmyOtsTef7DYbXPBxFR2
V+1dG4jjZ3q+yA9G/WxOfIwL8QeHvbwcNmq6srNDKEd+Uj4Tw3Xy9NqQvWKmdHKJt+Y5ZTIYh+6b
VGvT0Lar5NPCe8dAizJ99MMtqbEiNZGr+g645E/SAbY72nzL86vFm0bDIH+nOcoV6bwKVuJtNxGv
hSt5rV1RvbiAGLe+7aSQS4uj7SMLODG+ex831l/ulXQMRMA9xRUzNk8w7MhOPoFmfgq7zuAggDu+
Wce/HkVYZD3SqqbhjdfPyeMhGM5JOkAZXkGd8tdHW3H4565eyDcGP5fnxzXxfL4npfUk/RUmTJx/
DOekk6H4GCKHu+d8np8QIpThF0hnBsrhbTxSQZCPpO7ZgWekpXY71sOtCTp9Pk2Eyosbsd0wdPG5
0F8b3YoAtb0P+JH90WCe8I4IYFr7GLKdSVhJwuh8Ta/1Eoz3X9v8LPrUSpln2F4S1U9+Bl13EhXj
aQJqTwSqpy7LzUkBkhgutUSTVpSPRj75wt4M42ag6O0GfSM8AD4+qHixp3YgA5E0rSgpbRMZdrHr
8OBKKtHZ62OfIvyg82WE1rNqBH4Y64SLy54ty1AYMPLvSS6otge8FdHHqkbUq7Pzw8XcrSi8GL4U
TskLYBxTm33X/syDhH9Zu6HPY4PnLcNVbai7yUeExBcCd1vMoLHNjFSoGBoZc6Jx+mChRJEr06Hg
eXjYP2XZ1m0V6TgniingNiaKQHyQ05QE58q5SVbEeS3tGmZOKTsSwBKpD8LET33JFpcT8IkKuM0t
z199eBR/Z/OUdupilO7uVZz3biP2FIRW+6zMH86BxkSsgJBZPmcYTjyFEOg/nVexDDPlfim/01e5
TtjUClfCb8sSQRjn4zt+c+DQ+tAMapWxlkvb7BOPMzLIiIQoWV18NbIs7o5Drjird2uF3hAZq0Hf
AK7uEY9MUkgWELBmDVe9VHIz5gpRfaPeWE/Dti8oFUAQJno55Byy+E59nl+AYsgSocVYYz3ihxuQ
kqvKcJlDvW0xdXtNx9CQFAfmET2Z3Ty7LkgPGuYdMhfEiphueNjvheBEE3zHD+fsaVKAz2ODnQJn
GZWyOITHVonmy0LQ7cbp56fukvN0zn5u6iNcxofz7LHyiwwP4t9iYeOYHhacba+9r1J3z9Pwo5Zx
UU5WO3fjcFiaP+PHvu5VkqhI/cCHiy364134q+DW1JYZ0Kb+bY5nG0+i7ySHLsXdXBtsw435a62Z
OwklejugxXqIb1m/zXOC+ny3OOhbexiazXZviLeu2NB40jZ3o06t8YfhWWy4mk7WK2/rrCmn7YZg
bX7ARMNwddnpA9UkMfNHjzEbuxqEOkEKiovEy+h589/qyeLtpU4fcnJKuxwzep6VPTMIaWQ/Mxuj
P6LRGk+A/yN+yPCG0fwTS4v27+ag5oo3kmnfbNkFwsKd1A/onb0PWnxfMhCQ1uS5Z/vbupDHWnD/
lvtOXV16FApVrgoRh+dJyh7R2lk0AkqtT2NVf8V1yGKU0g9iJwu3ynVFpqpaYAJ52qfSU1Wn90i0
dAoqEy5zucBmUT0VxlK060F6VPXo5cCdY/gO2jlOaWi/742dpoiQfNzgbuHVeHYGsWEWvRZhJz+z
8PUibmDoGUorfBGLSaU/9d/DPMhEXjeDvxKdrZEHZP/ukBZiDkrfrdEKjcqIMGUbmyrzDOsbkApf
jR0kLU4Ew59zEDiTFpwA+CgMF3xvm3+3LWv1OlLU2Tx6gAuqOIfKPWnv8z0BuYwQmmr8na8PfXDl
Fys3LUQcn8UCAYZvKgQ2z2Q0j3lxDHYBnYrkwsWjmBkC8oNaDEwQhD6c0W6wLY5lYRLCfYsRktiC
gfMH6dy6GmpK8MwxhJE5pWAyhEbbsuPkWYBJLtO/XBPMR+7RjAd5y2Iu4F9L/YEdDA3wv3mgAEil
Va8/WkiHpHHGmwZADlFqOD2zOOmEkA7Xz/zzD+G3YXcoKHLb5q6BZHsudH/7hwiEDzt9x4UVCW2v
YLTcq++O2ENYgGXpu9R4WCB8Hhf5wEaoEXdPSPztR+pKg6EG3jQQFHxrYYQAxXIbCMuLKYBxmgy8
n6gm2MiCaSaLmTUq/m0iQjbtiftWNPw79K5HeNztbS3g7mL4SBvWcnOQxWEjz61bZnJQlJjVD6nP
YQDEiq4f5+GylFoyIRFRFCptPdPVXqyU5T/Md53JIcrC9oFHnLy7fjVgSVgPeOfMN9a8zdb+kiF6
RUhasmcxGUQt/hwlbG8o3b3inkT7MHYi73bF5g8RFwketX+ipZTXvdAacq2wdG8axEsrUx2JBUX2
CrZx64OHJe9Y/D7b99qphGbxLZhT+DiJcpasK1gG9qC4LqF3QsZSV3jKtMK7TO2X8kzum99EXjlc
peLsg/AOhCM3OJEGDibFlMrHMHyvEbgZ2dgpcvprABcqMxjsxlkJ6vv6vzwBXe8gkp5An1hwa5FJ
HCydFK5xjsyl85M3bzVjnzO7eZmRbUQTPAHNDNna6XOekNH3EbF5RvhM/lfGX7S/2z1z2xoI7ULh
b3t/5Kl+rfTG1AlCd0ZmaT6GfZz8YRmimYbcfE/sX5/AG+0BA/jpmDTtuI5RxoqGiiCenLyAXEwr
YqPta+Go6vq4EGGpVBlh0PsSo8O3hbXCf0rYUPoIWXf6Z7Ty0gks0zSSdvN7QjkWsTAnc91ezzdm
8ZYi0o3qEJEc6bZBdpXHRDwoenk+AnpIBk3ppgcSab/pi9DlCq58bZCDxbONvKuT3MCEupHjrnR7
XyHtYkYTSuCyLYayescIXKxsx9CeZr71Q9P5cgygKwDRE+zlSAcYIduKlBXwkBijUCR9nGkDmvav
9W22At/1OsBe7/1d+N2BB1C5lK+tMk3q6+J67Hyn9goPJmO5xxLcPUkW5ZrlKIeK5qLJWB9trkMk
rY7GL7dEkrh+xzak6IYkEhYaXfpV7Artn/xDw67lTLMsLafjG6l+F69ZHdI242rmuuSc/Lm27gdt
cRUpExHUi8GNdHsSz+RcovO+edOmma3GULML6GzHr+CxehC42lSuYmE8qX3Vd3RnTqUHQYnZqdv7
WsqrcLBqrBqqUh5sWxayY3VcEBCiEtUWVlO+v+XNuCHniNVy+EKrOJnT2w/Wq9JMqW2iGDs/456W
vvS0jVadSL0x8dx99RA7/g2zX82Z9ZaYLtW0xBD2TRv2pg+f/iRyAp0Z4j3T12K1S0IpltRebPaS
3vR4jJ0Uwr626UYMjtap4u+MsiqlXO8zgydz0i1vAwha3lERNcZ54a5/BSF2VyZK/stIaHnPx3XO
kRkx//EEnsegqxdNrPmrpvXBtaAvPp161G1m30KLMKhtukr5K823ZTiuitMDdziLZduc+iDxkXwe
Kdg3n2l4c40XELdymCURBEjVMspXyderCkjZt9JcR8vNJDMjXnjLySjftLphxiTFARbCzu1iYdLK
HV5fdSbjLpoeqnKAgQbVhQgF8MSCLTPSzP0Gx+W5jcgYuSf3QrRBhdDarBBbqvbjhUaGUm/n9biP
XdT0LivVGIoIP35NZC+aP1kowOCLmqkEEgDy1kg3BH6AAYaNTO55VYO23sIsRYQoMDr/eMFAc73n
S5rrwVgw0Ds9UDlS8otffdjg4q6IXqtdy2UpjaOaKC4BFyWHaFOXVUJ1N7CffvaSaDMaNrC16qNM
nf0q7NOZC9kPy2X+bUB1wujKxwMszNPhL8riqx7F5/HKw3vBEB/X4vq4Hlafk1uiyeZtNTgX8GdB
9bRLprHOF+phIW5brC7CLEyawSYIQ4z4KcZo9dy/dHhEHqlbg+dGyrtqPuBkce0u9hEujfA0W5Ls
xqdCtSHVLgHBqKcUqvlNd3NRhMpgRDzJMFKNYaRwz6KX3bDsx+pnvaqN3mj2z8T6jzKYKZhHYbyQ
sN7BW4v8Vj4K0vIf/Cdjn3UFWw3d6u/fzIYojAzlnat0GPa5oAEXXG8GLPMxODgSzNY5NkUmnw3p
Dak5Sj9EMy/s6PMvTyT5ym9Tm1H2O39R4P11qUrhg9Sbq7ulPUPll4lZGnXNPYequFGaMDRgX7ls
sqdnxEaoO66gk2TatCCNmUJ2WZnNQEhtUKN3UtIGJ4W/3/g/959jJ0kV2B47lJEpOme7GFxJGMPd
vVS5/gRGLBgu+TkstDDYs0CCtLKUjlSRllgH9yODPLtzYthDnECeIiRgWJcK5WN6P07jd5IF2elJ
ucLtkeWPx8DUIGBjAY1gf41rUrB+OsGzeWUci6Emxruw7InaHZ2kupKhyOGqQp27vLCqDKjiTQpi
PXgkoHkSeCA/JidvX5E4QHCjJxOrhsNEJZnCKGCt1vNeCZtuw338+Rmug++ayENjTBY9qV//k8ij
BjlB+168K1drIGY7n/H3wIop89pyNGYjJE4K/U0ViLqD/HejDERUP+quqQJNRC0ovFbQF9NSm+us
aoz6F0UpW8Bg+4YdKg8oiDAI7HQn4Gzu8q55EYk0RHZfcvMISBkiaJi59BQNt85Ufc4YW4l3oO2m
dk700o41PQP/luBIcbugP1TXCWjHWPUewl1I1m7mnhAsnVTDneSbY/9wa+sDBcUNuLOcDdO0ojly
nDVIM7b5biXVSxH96IZ3QLw/1cM5iDXR2l5fIgG9GVOrp1mEgWolQQdfsL3zr5GEo8NKGXiHzd5V
6XKJPuzMrYs2m6PDro/hh5SLcoT83Keesn1LrTBTc4QDLgwkaG7+hLoHBaz+jlxtxlkev61FD0Zw
1Oiml39j5XkC3NPaIuX5g9AjyuF3MLfcDmKklS0fYzlW8mI92nHeMSSf66qTvYcF1PsuRNGjcp9/
FjnoB3ZnBmj7RzET+22RVdAqplaBx8Ea0ZfibrvWon+xePiXpu+5eur7e6DFSlYx7W7g2XYcUfNS
mgGMARkkkNpLJf8e0is1cSsUAXStdo9Og4t7jZfbt6wSYVV4cHlQCgIclSEukr8e4PNcCaTci5i0
7ZRaOgz3XI0nN5SxQCa64zJRFw1BUkxQDfIyR6cVtCfaOv8zDs7o9QUwc5etuukS6OIHSA6665ap
fabJX9TItdeRtGhrsm0loNa7vMCkVHOWepCfINMVBnW1NM8oGglYcdXjxVvN6YEA3CQZviqlbW9m
E/fgYL8V0pP5n0HP1zKDRDXp0Wxja0NoqI7BMWEeQ7rcWTOZRxJI1RzpaZ0gHAQ8YvARMvjAAyx3
0KLfO7HczmnUyciJKJrIQZgJsjya3p2W6/nm2wDTHVRK16kbe69ffTdwq6eCo58LUH+JHI5Pg5VW
9r8+U6QE7LaPHgzd/NnrjvRlQ9GPjcIiHBdifThVcm793UPPbSh0vqy2mrsZYIrQejsHCAnHfYKw
plKnmmybDlydvsjDky6ACyyq6yHIm917VDv/G5JCayuPbD/vgamMrgNCMTcanZKiCub2ZB2BEXfo
fvUxsTsz3kZsrZT9F/FIoiU6odZJZbdwnu+MMJPKvP9A+xD0vHnTOiLcYap4Rsf37AHfeFOjJX14
ejH9p/mqd3L+u9570l5HggPUXNNE9+ToS9lnfrYNtIaO8Qf/moxH5/v4b+8er8cR6p7B9numiCvs
4ndAMj+Yng8QisIN9vqIyK6EktiJeKAmzZt7IO0aVk1IA4AjeYQSghUngriZPgLmmhHbJAhqxeeB
VsgbYSNfw9k88Zw6ZGIeScrt/oOyA5Y5t67RTaMhLEZTT0eP1Axv/7n0kvgiseDOWItbXA0EZj39
97hHVMnm4c4pmXjuw3XD5N7XsWL57b1dzlJT2522Re3GIZsU8+hJaV3ToaGqqoeXmtEc7cug6gbk
lZcjQJ1fB9w4IophiXrs57c3OPdEv71xtiZUIYe6P8L/BeC4fENX7C9MiFG+9aDoJHVQTqEuT1sS
NKXpFi/okn51W8lVCOGA0IrNyZuNQumVqCNpEAysEuaM4+Auc1NLM8sHDX36UpkhUcF8lu1kDZ2o
9mS00XYfpMRc0s3aGjPM5eJnRFcxVEmV/qdsKUH0Shtrkwmn/0BlkuqNzBxbrLb25WueX/7wbhyQ
bkyzfLok11fKDj34uKfrtZC1m/QqGqxUdzNAnwgC5jdUihRm0iSDgCAsSVCeE8XWBCklaTMQkD5e
K8sftrGHDUH7jSZUYgNtcgc2orUpukz2ExcdPKUJeBvX77+N1DkiQiLPDVeufq0+C1Em7SATMk5s
+Py50kJ+Ui206Wj/8gULmpYoG3PjYdcJvRkfmK91PlkKpR0HpeUlKWj6kwlrHVrazR5PKxAvsdGe
kXFTjicUHzpCfpufDevrqAr37Se97CCNpub23Ut1abKSAt40ZyIE4CQjvnQL4fdZwmRQFw1O/4p5
ESPJsGGygXdOTzbiLTWpcE+KrHsno+JExqVw02xyESfIGcIAOIdnjDImUgHwYTiAMi5FETZ1/chK
tgN0xznw8BbhAHnvhSK7BfR1VhTKiOJYsHv0gVYyKJbkR/6viyT5swrwIS0aRc/eAAT16bIdq1Zx
5adNuotRT/BNXs4Mko0s0hgy26MJdX8M5tT9VHUWclq79pf8kPeTBo3+aAhJetldS4FRRSSv2XIc
mpclxGIw+PgDiRY9Zm0o37BJyLr1oVmbBfpw6bcYxcYk/+Awkexmy4pbe1p0GNsaoKhZwR8dMaDq
E/11K924NoJSQPs10IiDJwr0kvzN5ddvw2JWyijxsc5hmwOaw0ogBhBjS5eob/1HIhAcndJxosji
C1OqNkJ+t8PCHXzXaFRSc3DltItq/E2F7AcWZmCXcsMpOCxcyWjDefa8xuu6f4ReEM+7kl8m6Jrb
4nNSZPpub8i2GdEeCuJYCYZvRnOZkirwUAcU0Y2RuTfVKXNKqD4EfQK4crgvAlUxglSXuBqi+EYd
2NzjGA+29UGhb06bEPEKs5jgpcMuG22kiHZXeFqHKmHtySfaqxbkt5aT4snHPzkewqmY92D38hoq
ijJSCd0vwCJ4HSks6rlyc+CcWmoRkSSGMy6tVI4f5D8YkSCtzo+QP7mWik+g4L36xtwp7K+7YRxl
ByxV9qa2j8+5STrATqhtxy2yH2x3p3AHV0TXQkKzKhgNa9PnRkv7JZ54VCSxcRiRc3W2AJpA2X3L
Ni7Lr6quZQiqlWEuG+IVY695r134djq0ND7VxEvFpV8hURpbFBI2cq5U8KPyiDmjF7iXba2ANxr+
9PnUO0AOoI2JZ1s0DZxBXc+UvIIahyaovblIYTkzW24vmVwSS9ICuAwAJnuuGyoNB/To800gGH6H
yjIL5QwCymUssYoGN8Rqpg7OOZkLN8hFt7/qXSaowMINUeecX2nugdAbl9VEHtgZlWwfbOu6SS4/
2tWqBxiCL3d0OwHqYVGWU9/4g0sXw5IKDgOy2yF1xyZqhAvYLZ+yaSxVl6QmrdIMdxRIfUmdtQlw
Y2SUlW4gZXT6SYHvpljb972QkZrJud3v7NCJv+hV/uc76h2AzVMs3H4RfnVb7HaXZtCefE1x2uK5
beHvPnV80yhJ9T/QxvAiPHpbuoOEumH5N0Cyp4s2SYm7cO0BIMM5u7EeKZm5YA5Cio3onmllBaKX
NcltuASVqUN2sI26dOtW3a/joKPaTUrztN1rTFkWA0J9bPyBGKaW6dzyJW5J3V63o5MQoPvK1gEv
u5fYcdxBLAwqXR2G0To7jgZoQrVSVWa9u75cVKMtwcx9kRF8JF7+4BFvK4lh2YBvbXnaBrpkakiC
T0591KULLzcmEFDk0ofSlwrR3Fp8Qwcv/h2cPvG21sVFP3Rbzebeze42dB1yTFdflU1fbAvqG2RU
rtVpk5143N0lwLj7HKM3geIrCzJsiGYqEkm5lIt+7d5aglg2zC1OYqVuwMRK6Y8JWDOG4FLij3hn
nTGKDiIX/Y6fjT+6iyhTBmZYLcfQEBLncvf6dEJlmXrWceHI8d5AGUsviUaMeUV0nrawGz54NdD9
8LWt5qdNF8K3RpN6F9CxpiWiwwKQzH01/qBuMkG5Y6fRL3mv7Eiv1IGMygWcNxnNFSJNyEg9z14S
Y5crr0erzFxCxgJtPz3JmufaGs2hs5w4KFLwaNRt4VvyHWeRult815qq6vz5/3Az7CrQtWksZbH9
YmsTdha6wtQ0LBcRS99C1oGA/mIdsrs8x/cQ/3wif/UvM9h73YPPlaYsVFU+dB/ypCY/jEkWRMQE
9rSf16NCw4RxbRRK1ilFGfWbcM3RqKiWkDMEanSeu8DYRZlXGtHmF4M8TEPGT+i1AFSWfFX049Et
GAtaryOgs6jk7B901OJ4t5bUP65Ki3psV0pj5LyAIwRqf17gRU3CRj+Zb2+v5KeW0pPHzZt9tsq+
tg8/YnOeHNTjjVK6T1JeUaod7CJht0xGi1Chm7IiflS6zTjjBWea3vB0OJH6PrUBaagJC5/YJLpt
ULi6VNtLUW032OKOhgHG3iEVjYp2DVtH5h6lXmZzfrsV3LmJRAJbHwAMqaShZQValfi5fF2kChxd
erPwEZFP2LNqveCc+grZaXsrdd+z3be7g21rNuuxRF65v3nqeNCtK4vwlZ4htI+7dOD/w17ni/kK
Q4fR/3IloZw5kcJ7sVtJ6Ht/h/IfKrulnWDkyXfbB9e45L5CPyBvLNag+MxgXSnuLnMRXzbybEed
dtEvzFUHg0qsuT0Iu5RaNMJB/FUnQoZJX4mi59YFgL/03q/Esj0W1oRGeJfPyd46mabetsHnZJHc
w/hdMWavXu3el0S8DO8PDel7dwe0P8xXceZZ4Aax5MJrD6qdKla1f+GK/r065owVga2cH6uu10YT
oRTaUAOM1SEw3ApOBZ0M+TLyqlO+LFs5HxagKm/KnIDSgaxluRGdEIuakFMXYni5ln+wwpcJ8p/f
YY2KDZMlRjqvlNcU5aXPZigNliKpamsmju3ubj3W6LnItNB2UAk8udibV5AXSTtHK/jFNH8afmHi
PUSKBXCnMK1geC9c04NUG2fwmT+TNnSu4ZXL0H7FgiwNspJXihmjWfwHGaeMCmTMdvEYjCVEsU39
d8vTsL1QU9doTQvNRS9Bg3+tgZuPBhJ3iI7B5/UHKuYlSmi4mmYgybu9IFrufTUDgND3E2BHU2vq
g/5rJpGHSU4gAmpWGSLqUkVRVMznKGG/8icaypfdLr5XGszrjo9MvOIPxS7uskBUZzDOHsVIzCHD
wgTpLyk8rEg8hNOQXAZHfXtP98qKItDfwW0I5G6pNxCDDPknawZJCCA/GyAc0qnSFx+sSUBm8ZGp
oQ7w5sw0IqG3fgiltIAy6b8uPgig7Y/0gKwDmLduYOIORYeLicn1PRLZ+K/C5ShIhK2m1U0clVlb
Pjb4G77ap8LxwO7GAcVNFEBSmgjVV/7czjZdFC4zhLCrmBZS0tg3aReyLfMsM5KWkP94e5MGwTJd
srIcIk6akNwidIC4IHau4IGJYRjY1axPM4iy8QUVs+k4lSwWNpbG8FpmAPIQhq/YdoKhO9e0nMMO
6repdD5/fzCyXEmpSpQoLuZsT0uBGI1K6W3CLrOV52W76F0zGCeEPPaVmZfI4+yMX+/AHxzbxJFp
e05EFVuYHC7EkS4ahPcVV310aI63FqNqFGBlxL8onZ+fMT0my1JTqTn60qaUanF5rXXZFM9LdkdW
+eubdE4TK3LakihygRbFA4SXFb+mqUavYmL8iuIWqHdgfij0S0wq5fDVFzZDmvRcGhVnIui8KgPm
sT53LKgX8jcl7qktjYlNd74M6LyamZJfdZFZk1e57thnP72nLSePr3WxMfg2WPE/HpjQza37J5vq
iej+q5gWZw9Fxm4wUlZ7QG/mM4r1dliPemBNouESmU+IYK2MXnQL8xu4PoP3ZxWz3E36wwKHeAIm
x9BRQaAp1eeon0EZPEN/ynjW/inLZ6GWfQ+ta0VsFEF/kYW//UJHtEPpajpuLc+O9D28rzU8aqgE
LCD2nOsDOjJSCFA5hD68f5SkNdZj7YLxLUckYfG3F9k6e1f7p7vZP4ZwAkBlpdwPS+XKDWbmkm/p
l5KSR4Hs6tEyHYcN81jl6f2tWgjil/2QlLRFANMVS7mTcgvtGHiCAwNgoHBy83W37/AGLBglO5YL
NO+VaNPNs6iYz02xaluUKeg6vgV/UHrvDoDnBU3reTj7vIuzEfXwg/vesppZPHMG3TRiDIMawEiB
Ni2MbeKMpmzIkjjwC/KqLoh84B9wxfZsAghn0panWwKKX7AIuVFxaIFacWWBHkWZ2OqJ7Ez9aLhe
hq5sMG+/OVBftj8V8GdkPeuYf4t2rjoEeuQB/i+yMKPeQdD1lvvmXLP6d+75SqkzIcGUDz9CH8ms
7Co2mlTx0aA4pmlLw/qb0+lSdhHj9fOiLYsPYSdLEEFgelX3GX0/whyknYat7D/sQ84qJvRWTBDC
e4XbRvlRLH8cGNFqBb2Cm2j5n40Jx5/mkofnQukXsRsvcEkcOHHzNGFtnKdtYlDvBT/mcLBOf4Ob
F0O3MtTCclvMQaCIt+N8ybJx2vKNraflpNDVi3s/DV7okOt4f1XEYHxpqOT/qIlGh5Pj6YuWQX7i
YJTpiD1KZd7u0ZgvTBYK+Vtn9/vVwvvyP6lJcjwUyfnH9ePN6+M/+zcx1K6HZi57zhLa4WiQ3SeN
ZM7tpX0yP4j3Titaa1ZUmxIlp1znzY5QfmbwRpKa8dk4Uzjwf04uXnwsmZOLJSz9ktoya6y4nKJH
gjl4jU5A2wCq6Uz3yp+mJImHJq7mSMlGCiCzlrcqiOXrXWcy8z/MRspHZ46ur6UNFgHkJRwt/Bip
/gktCeGa0YjnIZIItNHktOfbgGLY8bv8SGbOKlVQPXzr02ibQH6HojBTg2K5Av2wJWiYeZorWL9k
CKjZjW4ftuIhWfIqDyU5FZwWjffpAzmFiq7suYpNMvSDHAastwCg4ZH0Wald2kuk51SeLYnrrDWl
4gRflTkxiAVK6QO+p95udEGftg7osXj9sRu56jB1wcKgoeBmVSPODOtuogGfUgFSvcj49IzXWBKq
A8jalb/rFZNYuOxtMiwAjdyX1ALbBC2E5xRM8+fCXDB4nh2d0N1u82G+zu9vPHh/yBQe55L/L2s2
BE3ZYNTr28bT3Mj7RZMsMwamfEuDobF4BydEk3E+BdEe9V9PWBJgWVm6nGPhOrXVGxMApGwu29VO
tMi0HLEAbC+WkGVuKJJ4CfnLufZkm/0tYHBRK3U0IxuNUeDDaOItLIyPgXP0GkOfMpvQ4k1oKlOz
tmghA6fJRwEZYfZD4VHt6IcQkBKsKzoxXWtAJQ10g7+rstsVCmWvGHOjEx1Mv88epC9BiCW/Wrl2
yLB3PxsYrIWT8zcpzhtvdtO0Tnq2O0LDxoUnPQI5LifgMjWdRaBBtqn+WX35sKIDYqRpGaiz1m50
0yDgGO7azS6sqyvE14yG7RWCQa2GrYjxafW+d+r/gaQ9SYFk5DZ931MQSgPgxfISphhzWMKyq1Q9
cewuYvm55c9yJ+U8KAaQ1IVOGFtLZeOu26M4pxInoufiBZCLBM3KZ4YLVrzNcHwYDnXvLtw2x3p9
RMPXICQJn8YbM8e9V6Rd/WA0I6EBgPRRITT6kSq+LIkiR08Eb0GgTy4Hfe2hi0Gtw3GpE9qUL8f9
ugZMJspBlGwHg2bJ//jLQlRnsSUxqKQqN55ia57YT5yhmPjcqnDT6meNsNprtKgOoFIEwCwFPpAM
hGeGiAZVh+iE4+pED/+342Xa+j3FH7Fd3So7jIY0iJ5Frgj52ZQllEUrFxykf6N5+9C557VsZmJk
9KZK+9XYp23nxYiuofXz97eg+PtGqmfgWoqyWJEY6RbEWuhHCX5agjN7Fa1pgie3ZyEoQIGkAX3A
WeE+MzS3HzbPVz90DWUcfzk/D+JuYJKEh4pz/o9tjn58sOzrCiQJp04luaSn9A2trRtM8HkldcDe
Fig0R2kubogJdleG9Yw93NKjuSWJH/dkx+TTK4B/ZOG9ZlqhTYoZIdk7NAaaQnZCj75FZNjrZS86
1nuLW+4tKbJgVrNPUqojN0Zr2NbOE2CyetuL3pxG/OqnT18ms4tSXK2I55PQ+I/og3h36ZHR29FL
qRxlaHjGiClBcpmRbwLtTjuHokSCbNSPHVnNb4O8G5nF/E+Bt9U14364cO4UlNNjE84dknjp+Xwq
PPXu0G/GuSTG4GblzLY0NrNhm2PN+xt7wkMeOqygIWT5gCxNo3ZoisSwuPMvBFBfTUxdh0bLjMTL
gBtY1kZwrTRLpiCVo//jlRVT7T1N1tfChW5eMJDbUhrLgBU2fjp2K40LDrPALTsUlSSivrtHG1BN
oHElwLqx0Uo1CtXqgs/YnWY4LZYbwvBxtAXE50ZZ7RhzFLdXoh/7N5QWDFRKJmpnFWkYK6Y63D6x
m4pOcztt9kaTZlDK0lEKD+iZxQkq+1FE8XnvqqDu18qMdX1XOqGJZxl8X511ekuWGvcCuM0Xy7Nv
oSDpMVIbyMJcv7Ow0dx9P+pRFMNraWPUBz3Slu9v6lJus2T2CC/OIzgujiihDpcqOtZ6Ij/IC8Rx
NsczvckmuC5vMctzeJ7mQBRFrSKUuurwNY8enTuTv0rOPSDJxSwAwEVfKU82OH3xUUMSWNt/LnbX
7SBJk0tmWKU0/LvdB6TLYWhwUqjYa16n57fjFJR2wPb4TxJiboiUNr4mlVWa2XcTQ6cthBEsI9P1
DdME0wI+UCQi4OUTRqd5HC76nNBxQQVoeTP4fx9PeLf5rQ+HK1I6B4gj5tJXilSLfYaOGBSxWeVD
L57Di8sDawUFCy5UyHHT5HG3nKcDB3XvijFlnxW9YUXtDnJVTUvHzcPwhuxnqq0/OeOVYk6vlRrP
kAQI0Ob4Hp4hR6wZz4VziiooomnhROFUhjdGd3rB4lm9yV2lqTFAycTHeQCVDCFgG9gseVPpaQcX
GgYcyYS+5CcO8xr3MhaxNU4TUiNgt2xSbT2PGwVfcg9NOFO1rU7hRfa/jU00R7GYLu9ekhzwiXaV
tRn/Z+wL26cpOc5rOhOyE5208V1z0eJi6XYf0k2TwkGJRnUcpIHthp5O+ZHyK5JVt6Ot2VTTPjhk
lNTdiZOEJjbVl7JcGU5rNa8+l4WRCGuTp+Cl3emH6bOduoDEz5E0qjmvdMgpRZwQzmIPCpq6s1Y3
DN3PgZROIiK75HrAemLv2ORiQXmSI0+aZDv3yZ5L+UlJMC7VFmCyLNHMOVqVEhT8dMKVU9KQT1mz
stZq2w5v4tBr3nu4B73twU/GKMSRYdKwS/h/xALDZ3fkdueHLtNWFbpsgnJXTWUDKIdBxGZq0TW8
dPe8XnvWP+lDanFes39A4SYitiTpQdfcf6DMizwbTFfnG5SmHsx7Y8oMN7iQfWWAFGXIy92a9J1P
svqaKLzdkwUptBIxJzsBGAR5KfrOLuhds0eWDFKTo6u0un1hzcyUOgNQAuk/TjnjWPxxu5gj72zl
REaS7hE/597LeY9NbCPXt0UuQp8Gl6WR6UZppg8ponyyBcy1RM5fhBZsVnP3yuR0swctOyvtTKyG
EfFwiqoksGmw8poDsSNeTxHKaHTDGTab7XZ9Wwg8EerGuU7ZxNhFW1ERI+qNA34zNMyvAsyHwYSk
h8arLuzikyqQPuR8EswF8ERTUvoxhR933HpvNJi3pHwmZ6SPwAJjSHPqMND5mkL/UurWbwXk8rZY
VvVLt+WgNeiRqUuoRs46LeJvVMJfrMw9E7vvQ6ommCc0lw6TToqIfM422p1/xE5HN+nzmwELrQ3W
nd2PRsiatVwjTT8JwxjFEte+rHh/wEGo8st5McOBfDnHoyjDXVu0ZdKPI6o4j7Lh1fFwLhFXNoyb
Sxj4VCztbpwmVJ2IBdfz1Qu0uYpgLaGsQ1K6/PwClA9mzuR+j1EKoCGw6dv1APJ04vjg+/LMK41v
SRpKgMZFR/T14XNPurpFt54mBJLP9VKzRtqCrRy/2hBN0ZZYhTBTKWs2MsBrGwf28UqElLLnRRtK
qPbPpmQ96R0aIAxHM2k8qmHP43L0X5jSnQ1M+V4crjfUpszibktEXbINOJ1B3RuZyNXMAU0B/gUF
tLCuxtfygXGI2i0JWmoJE/BB6XWFaVLrm+TVj0F/gfPTBt2TDBvLpN4YU9zEM1Bf7XY4ypY1K2Yr
fw/Fp8RXoKzlvb0W+peCb/TpDIXpx0hjqHAgtNV+Fhn4SCe9RI35toCxcHbQ0XOMyYKhxsFZVaUI
E8Fjj+DucUaqA1IXHECrA8p9EBvbciAKgLmcAGpip3EiMVeBFNasopu8VFIheLhHuT+/2hoXIEaZ
raEraAO3IGzHZNcc7n2ysPetN4jxrrFHa3oPcg4Kow82rQe4C0p57Q8VTVhgeadDlhjv6M0epTxj
WqmTYeoa6fgNsm5Uc2qSeiYnKcV8JXulWHnw+PVqAX+3d5UghvbgwtxM2CpCke50DS2fksUWp5Wa
L1UXPZJ+p/0+HL89kyKMufQ2hg6HmhugqPCHZtB2F2NnHuA68/AcMXsRKxo5IBdQPNR0/lVSbETU
vxRyBMAC6nhQa4bGM9ElkeqYvU2xLh2XXIUaIXztuKCgwN+5X4SyciTH9ZNmLRY64SPBCrH8UZ4a
8Ba/RopFsF81NhzK0hVVBUQb9jnVOU+dBS+TpcBOBdcVL+w8JBkye15eFsszJ3XPACI3wrtE7dfF
BmCAd5H8jd3VzvSsav55qkuyus0x2JChEN1hV714Fhi8bWZ9f0jcHIT0dEGcCp+njMcH48Ufqj9M
qptGuYxd/zSX5zfd9kHQkglBhATzmspv56yakxhVtzl1Tx0J+4luQMqCo0d4d9A3oRrtzytKmFpA
dP/fVb10mTbBA9fpGdGD3fuTOIb+dREznjGn60GdoCpPJAs7vipjYXeWxSMgbdlK5UmSe4oogub3
1ob+B/+XU/IQYubgiAnRPEVlCi5ufjdS4WBOtiG28mKfO7FCivpl+q3GYAmNp9qvZggIuz95hPgU
jVWyKQZTGgUYuybVpHqf+pTdhlbu00gvmYg7VC++4imyeVkVgXnwccELCc3T+ZSUzaSnuSC/yNDe
JnfGwn0F3oOWNsNF1NdDai2JjAzBDQObGvMoRitK0FcwEU2qZpfWmyi/ZlDAc3GJx2dNj/FFmIHz
BQbJAz1Qx3hzn/XR+Pgiur8XxzxKEdmZ24Sl2/7GKVySgdlWVu/cUmZdpkpxbZmQhksdLDasIn/5
xX2x7/9zihPKMYDAQ0FzQ04HQ/P14wBLhYZjkpuGnYH71LEYPVhXXoBlq+lJ+v2P1+O7fsuckN8Q
5uHWgOWSD0RoFwB3GKv4xb+RQGNtJy3fI3UUXK0QvB/77GYGm2MKaSZ5J527ZLfAp4o2rYYdUwHT
6H4Pax46mOFyLBy9oXQx+71y664ZBTjfpxYYAA8IBRl61ptASnQpKxNJc5VebkgwkLcY8YV6+fZJ
YHxCc7bwnu/3UQon1cncr4+CP2oIgy5EPlurXja+DmjdztCSZz02bFs/kBxFNniqC4H0YV+2SsoD
8dh5xh5XM+oPCCn2YIF+LWPmexutAwSStN6WnkQc4cqLG50KGQhNolPbcZC3H4dft+x3O5EmmHxZ
VwzWuZOzQWq46vaSy30/blTM61N6vatDPQMyt/yZWW10gGHFMFfSGKg6hZw65gAcTksV9Hzss2BL
XaMMUbAPFXB3Z+Wtx/4F5HdDAHaaQC5oZbCwSbxbEXGVnI4a+mi59lJk/fbVVoFxRWoHqPZHCiAW
nQsPySRXuadBh//oWielNN+LZ3OIhzwoxzSumfK+/PDt3RQMD6RDxtDz8TYyPSYXymuc3sjK0Att
sFZJQYcMXd4U1v0AwC5C3cbd8cobCKC+gG0zSFziU+AZOrIDrUo9kTyGBUHMP0nh+fTZd+JdJGkh
fnb3ZfG2Ns/0mbNKtEpthhm+MMXWwmszo0S9WMMsnmoIqwS4Dxotc1CNDwddRQJHsweKiWbbWCCG
nP77Ri9PGEM3Zs3Wm7VCpSvh/tc8iKh/dYrKaDd2selrenJaSrZ4j1/M85h593M7o2A0W6PASWV7
1accRloXTccrYaspMGQXTtTnr50Qbuy6vlhF8Xq/HPkZ2S4G4qukKKoLebgFDQKDc5CtK8/f7MoE
BjPVI00AwrS9TL7D4EzqIfjfY2i3nX1uIwslfZhBQNgKs+9TPrnAK/6+vCUwyblRoJbBVcq7UtEP
wskoNu+xZpW6ISZ6/4f4Ikzags1ZCcTgvfCLcjjMA/46KQa7rs7+jxBOsCFVWl9H8dZziVlTSKPu
aGNN/o7t79n5QdggNaIFVUTqDzaEM9ZbLRE9nLbC9CQdcfq/cFbD8+u/0e/OAb+fu/1Q2vjpqPRJ
zkEtaiAxmXaNRbURUaZQUaafJXwYcGdxtSiacodZxrmEV0wCewmJe6nvSZPZpMIAFSsHGW8XYXeT
7dbyp/ox1aOBuUM610c/lE3KqVOcgEfkTC3uGQgm1KRVJYw/YbzRl6ALwd7+hZO+DmZy+6YrV/5a
saBNV5t3NqWXHq9BxOqh27Ehlhj0DvLgL3TacF2U2BsYks3GfKwzgVXfRMGKj559SOIxgON+2COo
AXmItTPD6i44QDHDVpPXRnbBTxp4oSVmLa/WFOsFJ7ep2itfZ0onYTfdm7V7jsL3/PKE86NYuTcm
350eb9CCSc5/SFxgUEOu2DGiOkmf1Pa4Ckz4crH53IgTAKrSpMTmdP2Fi22DU4LOkkALC/AEL1N5
Q7YI2GQglDKIN7MrjAknD2Ty5tycXljWJSbv7blV5n6BneXyJuf/F35BNGVF77R8VBt/0GHyp0WH
lKgEC0Trzmciu44SO98tuEIsfBp3qwltnofX+ts6+I8uxh6D5wMifhN0J34QZTQ87IMKVBQUZqGM
AwyXE+7D0K1zRxUV/E6wSFuwZfd1OAliKsrSexjdhDr6MxzCZTvnp4UoWnWSc0pjMhhJWbxaVlbP
GEuDh20akXe+B0gxjphfyoX5Rs9fDuclxzFsmGmyXy7yFtS/s/lw3UgTEOPA3goT/nhm7VRT9Em8
jZlPkfTY4K90Jpske49uSliKwILgPTdb6sis2woco2zzhCc0aBC1zzhAShwmfNY+1PMeBJbO3GZv
7yZaDk0qhzTjhnVJTvwDXenpHHsyF6BDV1rHWtQxs0ecdLEJl/zwnjvvabAonSjr8ONhv0HEChQV
LeaSKwh+cDU437FYNywIBhkbciITY6u2uGhzP8VI5TPpjeu7dF/zOiTL/s1GDV5U8nmgLdHB+vSd
GUGQCRpN45LcZ4qWKj9tz0tsLBSPDQx14FuEKm0a+Ary0FY5rDJcRwTSbZjDg847U3/e3uXavuH9
7cKdreJErJaOl5W8nEV8ZvvZWsQg3ICEUK38XhGZU3BAksqLoTe1AphorymONXsNtti7NS1xM1Kw
HH8SFpkeHMdqFQtM6OENZFIuhGtUx1OvF7hs5Zz4DY4zif2dVgHB/z+GRbrD+jbr8yRznZiwa0Ek
bgfZGFXXQmP88uEjYRtQ/DxdiXTpfX9llxcfAx32jzYSDkqXIl8Sx63bUAv6k2D9nztB6urufpLw
5v9mIeXMKaduzodbi8tvP5eW1vrO2hrNZZLVOfbw0D3l6YoguPjiOudeNDZBK0NRla3tyAxlSMwy
RwXF2XU1SOz5MNO445A+lyX2sZZgElUb28nua9+69d57Qrk2buOTqqxiZwFE2nVgbH1q0lpuG80e
87AkwG0BTIiUTVwL3zbFhPf8YO38nZLx+1YWgw44vC0K8UZR9PylFRX75Okq5TfG+rX0e51d3ZMT
19XTzXiuiLSSy//8bfVJlJfU79H35WkfRHBZN9XileQc0GuSf5kuz9LUzJR7U+og8iciuREugm5z
Sz2DLeeABBFrWChuOWDNBmjSUijAwXjF/4uifEROReCbdp6VCzAdiNgAmkNL9WIQVMUv7H9yGsiO
GjDrs7wTaZVbqwwY4T3YCgEvUL+HMBIMi1j05PHVjK0mIFsrI0LsqtzAGEYxy73R5FGMADXHoywm
ZtwnDT9t2xYQvx0zGJZLbJS5owGqudrgXFNo3/nbo9n+9QGiDF68vRlktWveE9s4nxm8lGPpSP+9
uF6dMK/rBAIN+3PO26GJMQsTfL/hj+h573aFK8hT2An5cXLXkcFStjEWr8mRVwhdLy6YqDjw+CXu
MqnQ6FzRZVuA2tFnUgKBbeQhsq7AIXlEgJpdS1vwsqzbnOmdALBN290wZ5YmOV+hVhUsps79bdlk
Kn9x4zSgO24PpZ/leduz5mUa0kgGD2gjMJUGqdkorASWjWfu0fgWr338vLHxbzIyAbxCZ+vz5lY1
zWRw7rW0S3DqZLYpcc8rBaQxuRkyEx9ih6WoU56JBx5zHQDSqk5dbncRXU6shx1tzI64ug1fXMtB
l4hSlo0zJFHJQ4BB6pRnHeigxMS856P69LJlB76YB4ridkXNz/ZjmXylE/7f4dgqJpmKmdoG1qlJ
nYNd0LBRmBzQtLO/m4QxG7BX9p594Vpg1RqjN/49Ukiecn83hhT7AzfPck6UAU41dFVs0dE7Fffn
28iY6VVkHz+8+eC6SpitO3vzXJV6ZyMl33AjTtcq/7ZH3fRkucpTK5X+HIaVIZUeKK8jQ376J1CZ
SckDbkjZwj0lY2wqJOoPCXmLZ9pvKhIuuxBOV3TdezQluV0sWCExmLQEuW6DUVCTK5eS6mZroiBX
2GA6QjjEBt9laNgJzIhL1PWv6VxIqga8ua+D5UyeE0DJvHaUbWrAlqwjkBI46eZ773rbhKGNx1ZM
pcXjo887zOOBUwtae61WryPhEAT4ZLjY3wCwML0ozueAe1PNjU8qZe7HSi95CTgVVmF9RKO6nx9z
9/x9RbQRBg7bkewuEaCOgmTKzW308L3ylQmLt2xUDk9nch96ElEm5OcRilXF8tNw0jDupAxbM3zG
jKF8T5IgJMHzAlYWDmq/jL4CO49jdX36HGwNWkj5F2hnu1sArMKoTpeJ3Lk0Tz8V44PqVEhiG25B
Aij6ix8MYccbOho0yFPkNNVYdRx4mNOJKNfjd860GSu0tmBgNloKOau0wviaBXoo1XvpyZpyNuVM
/THPBZEV6DZoXTkt//UJOkVwP10jXO2aoGOFyCPv2nBDO/pGaBM9/iw23edXL8SD3SKTqTepw4Hm
VxslX8X3z+xr0zQJiLkb3hFxbyoV4BLy8EUGJX49BDckCNdjVvd1fWnXJBZAKGiVUfXTv/Ld3Gi0
XzJIfWYzZr6LjSsF2P+4QHjf4C3/KwmtDvvDnZxHTDCotnx/Gu1WbKJXgVm8pJqsb1oHtqyLBCQt
+k8ZcUjyNciSmOl29ZGkWJaeeMr8CpNjbuQR4XjfilPLnnvinyN5jmwz5o/bvTgsVF5A5mOgqL7A
r/8UULIlK80F0cwcgJ+b9ZOc66mheXs3q8fCdJ32Al4zAhg4DSi7FLHu2BElEPj+yYVuiqSIh97h
DDjrt6Rno3qtgAQh20Ssxuvs++QbvhewSRQLGdi0Fe9YvhTbZ3P6U4DrXi5g4o9fOqi5jsO5KoWw
ngGpqtmjSqm9+iPB6+rqF4Ae7QJrQKcfmuQK5S6oszXrJsChDbIZbVy7e8TBx4qsNpASJ9uqwA62
kHIfl0RRUGiyzt5fM6mAH5gsS5WO/VaMAsTr0tXkOhqmFzcLZBEAy5qEMjfRHeutPlsUd8nr4JP/
U+GcnGFPJVqMWZXMHmPUJgIMi36iy/X8BLyjUgqcPaWmRdB+MHdz/t9TqkZjPzsoxuXdh9C4c+z5
WmCqDSlc8ciwUK5+0/RyIhsGO9QzyTsHg33iwH/ZQ/NSNk3r5KM8sSLykaN1n35DvsWkBW/ulF3+
+jTqcYyf9V3zW4bv/YGcesYCvMiVJ4Ha5Ee9CPkIJwnZtOdMizDq2NcnCwuq318EU58Hd5nC4O+0
8kh/kiEDDwKF8rs+e8w5c9yLjJxiznAiQmVznPy73JQikRvwY1w+bI+V/lYIPyrdfGtGjER0Upkw
hfN8BJ+Xnxf3HABUKGrymGEUJ1K3LADqxpZa9/poGIMQh7s51WEb29jmGs5mEtgxaneM6x0GiIED
J0aFpZ54VVat1IvnXNJimOKEzl6vremTK0Oaj2mskeawxcqP6EJA2xrIyle7XOqpyNydkZ3/5Zr3
z5RDShKQrvOWNYG10I7aDP7Ere6kwT5SAU1gEHiqwB3sw0lHZ9tWixDtEWRNQloQ1UdfVWdSPpz2
s1Ni/fB8XXg3s4HkR8INTOSXGT+J3kmfny1dMhjDR9L8eiDsSJtJR8Ep4outwbdcUsEvbcQ0kMU2
ZAkVaPB4L/neFjSXhsYyH0E5lQw+dlXTNleo8EXXH0UeUUPtWLq9edWNOeCcvzzJy4DBE0Gz8iPe
oC4ccGTnR8BLaO83aSWMfMvb8ifR5BWbssTaLSSwn0SlmbEm5531meE2RUHQCfBpYqaQB0DqoO7M
L60tFIcfUYdSj3BEUKXmrZJn43CrGRZWYn5w8LDfYO50y41fo82L6BmYmBqQbLnYf1JwHQRALgjY
3gppuANA7fmuhuypzq63+pJtye5VD9SwR9ubD2/yvFOEr4My8gAIQDrgCOIWh0Wn1vujrLmO3Ddp
FnSRxygF5f/Da6sn/qaffksm2LCcyFkRY8H5LQDXv2WouNFpHHa8l90jCTMCfJQXAxyDp8eUNkLL
jj996DuE3kGkleBk2g5DDWx4Q4XbXwRVjlKqhfUCsG5K5yxcivVfSsUU8goYJsDhp/rSn8rNTxCN
mSSHy4+NDvCGU40KfbYLlH6U6QjCvyo5PALRFxD+yFTRaAtK678Mym9FdfpBBT1TqtEga1Ctiou2
n2ElhYeMbVwqYy3/b0gDZH98qec/B13Zg+h3Z884l/mFB8qlqD/7KKKM0Bh8CLSWnnrlQb3jnMEL
++S79iMznFB2pCiKZHYEUbVtfj9HHRs6BhrXnD7+3HzkSL+6noa44WcjtwDuxqDX05tysZoZ5V3T
DqA+hEtwzZfpO9TAccUVQ/Y90Jx5sKWOiG3Z/laYZxvxu6KNE8rmOa7aKj8nhXdTiuM2hgOmtrbX
PS0EihWjlUbSyLqol9/tkdMRGjeXMfyAxahqtKtQLVMxOYSoN9hDXNvVZPiFky0BMTj6vA/6zBJB
93i5Un/E27ZtOljYPBf2JdL0ZFwvGcGSD3oV8LJHp1wA/o0HG7NoaVG6NCQW7grYW03M94nZHQOH
p5oBpSznITaPujZNtCl420jV8yw4YTZdHIRnblbT7RZLjJ08GPZ5yXUgppZvL3krHQUAaLZiOg5x
XRwiWxUbR6Baa5goaYTN7zKeol2fYZrc2FqN1U+bvJ2CeNxbIh/4QJ75jyERoE+2yg5yIWaMNEKK
7PwknrwTvKKf0VDmeqtB1zQhXcL1unBaEGdfBLgxeA8enjZsO/1H+FHFSmAPY3Cd6mnFYqrmtZrA
b3OplSVolnsPa8n7U11DAa1LadJ3Z0CZtz2OI2NgxywLODWy9LPYkrmUPl7IRJUiVRSFGheuyaZi
KZZiHq/77Ry6yJf7sOmN9X8VjSJ4DnWh2jsiJb3n9TOYfaiyJL8y3CrXqO2ASjOW79N/G4lFhzoi
1+an17O0cPnRtCwo2J2zLUzk2OrYFisJkSWtGe194PnO5B7SCEnkzwo9ad7+sK4RHLxqS1n/jf34
egoDHPL+dd+fNNnQk0vv82YkX2uTBm8pT2RdPFoW/a/GtP18saeqPns30GZ1LemJDP+R2BwK1bkf
sDQD7SLb0q70aWVBB9nX8oWRkYk7YEiz+oXgq/Fc8fERyRj03oOJuUeMj7mFvllroRTfrKnVFELS
Vf5DiszQiS4LGBF1bayswAn7fOYfgQ70YthBBbAZuBu8k0NjcTUU5hHtwUQaBSmuneV749xz5S8W
yYJ8HqpVbd5TeTvAcwInUtI8SS3km1dnK7Ea6OA3fCQxLys07+vYKe2IVh7qR1EdZTmwFkm8c2bX
b1PLlL3skTnjUB7bcF0p7W1ySkQv4sSIYSU5KkJ818lFZ6/rr5UWWWZ58ho3U8ICYtz5naKcWB2N
4e1aC9jNcz1D4Afll3ge6eLqvO43q0eVFeE4JbrzBGqEb1r/iUghBsu7YhaWcrG3EnzwRGGoxdO+
QNbvu9K8SPCml/WmY47b5HLPgZemF1O4+sSmykcsD7p8oP2yW2+ZOSzqGrb1Yi2LWaJAxTdZAzF0
SzMMYvAO4/tOwQxOcB/qiDxmnhHDkbI7Byd6KnENRCy2zb04eFQ5zFaLZCUuALVrxsJD4QMXn3RF
hacytj9vyyMGcIhOn36KfFEKk3Ff89L3YXrsdkFkseKwEn81lEz81SSFjcSTdPp5JncfGKuI+d9e
1r4wzaB+8qd9pouJch65Fqt4eX7q6hoCZp2TYHRyvG0d1vo2nWIQu6kVKn61quRwxeMJzaXP9aHp
x4EO7xMl2V1YTNah40RKPzTV3QIaZeBnCh1k/gqhWjpilA6ARAa0zOFmUcPigbTfDXs66VNi61ul
q3Pu8JVITmu63OGw6Rc2JgufwCAjRaUNfIyMV+3efdHXyqRzyomcP2cdGEUJhBdEZ5dmIuG+ycIn
JcnKFSxK5RVS4yxSIPo0j8GHy3cuQ84uqtraRbvGH+MR1ugBnZAjC3Zk+qoVxwQWUcOS4WuyAIUr
VEsUijMp8pmPgdtqncQBgGNOlFRMQq522kxNEWuBtTbU15MoCr5nKldfdJuUksURu1Ucxk1+2z2W
jm1Rbe2ccV37794RW+zqLMQnOsCdkmqt91STFEP8fmO9YjZ1yvW8hDKdrUZaxIBlDpucGvWX5DuK
NUVscooT3uRFYCrF50UAqgb03wgnI7B85OXmc9CpgnkRFHXI/UmR3pR4KeRMFidataWotXcy+Ust
FL4bWboHAR2ejPDqWNRbWPr8iyXEoV/Gkp6bMbXHCLClqccrFUKD3TWB7lD/iwo0TtnxoyxRGcqH
ppvOo5lqFMLHlEZymobaJXKrWzeROdg+/i8xZVuneRvVMpWqa+Pobt5BYlB2nqW1ky+AsOMdLMla
ap5V3Lk3QBube8cVsVWjmlFPmZGzlnC2FAECDmnoeKzJvgcv2e4JvlkU9u/9qkLJeSd6g7oZdlZB
AhqM2Hry8Kls/x+J1FWvS9GQsoXn7fVewUGRRmjkYHYyBqKiilRpDZj2v/VRMblTq+l/GZ0+BE6W
ry0/m5tvvNc4xMAQCAG66uYOFV4G8B3DgQjiXYwtfwcFpsQGO2Rup+I0Xz15FoyILpa/ThpuA8Sw
n7U5InoXEQWzzi41aazks/uxJD1Klx0n/gIbkLUn7djkd/n88REbyzJJccqiclTSpM3cz9Gknw+j
UEpgKy0uqbah3Nr5pVQ+YmyaY8i3IPWTBvnxuhYXSFYMMoUlJn7ApTqhJs8jkbtlobAE5thQIrNp
CWTz0VW+DjEvwYItUhYtKOlzX1LhcNkDG7loYS1mCWn7brnAOsitJPwY7RG6jWje9EE6M+biqtVU
/mN+quiUIvXTTmyU2pSpYj0vhUFaunsQ8g+duMpBeFjbdbC3pqmuD3gUiC3GZ8tMOu8ua7cCl0ZK
iM54/e+eVUpgFG1hy44VkI4UAiXJwoShU1LAGXTIf2eSirsYsLB29n8CJFZUmTtZN8sokI6tbGCm
RPqzWnnH3nk8xnMoBgIciqy8KAH0XArdnL67Yh9w8r9hBTjiGS72TxU6G2x9fPPinmvK4yS1xrYw
0BNrbdSkhtEdkFcph4EA19Ky4xLD+agHqpO14m1ccL/FFW49I3INgnuey3x2fRrPMlnnfUwdKNjF
XW6WcFSKW94QdfmEssPGuxFucLLtkihWGvlZdmemFpoUOfFvX7mkJmNhlN785+TbEz9BA0w55yRC
yqK1MVdqeYgcZ3cZQCkBlTCol8hFU8ZuCJSjF9VntT+N5umtjRmuDk9KRlOqUySwrqZkKLerMnZZ
1lUq1/0hoE+ghaQJp2PSqyyvkIy3bncmt5HphAMfvJ5dkIsXSLcDuvTN1p4nFtnlfB5d0a6WQGhy
5k9FKk5hs4NC7QvrqDwU0R1ONzfemU6U9FKJJ33LV9YR8S9N6DSN1KRP+C9llJv2Hd/k6KQ0k3o5
6/kIXzYqOw2mESuiplwvFJ3ZdczbIkoFDvmMgcr8LQjIGK86tUcN0AIN+keOnioyqQaRGevlICHc
mJDdeUKx7X6mY11YSKdUpHrJAGP5dR3xyUdHo2DwbyLIU65+7PJzotyOlLeq/DnsjIAqYWsmsvr9
evEIzGUfNn1UhyumQEFaB5HWf33Grm/ViEYOrzHJqkx7A7sObKq2Y+WSNdJ3K6vW+R7KHn2J/tBC
BJ4W9ZS3+s3UOv3lSI+NpQJWSz+7jTQlLBilYBobpnoHYQ4RLLkrzSSHW+3+ahZQGSj0bDUniDFH
UbUfSyY9TogszfzFjnkMzprioDxysqjraI44CAhWczwkKDbCzAt3uYz0KrdXXzxjuvLSbVW8/AzL
a2u7IlTEeRVlt72b7O1JNZai8byXOlHPIBz85MMBITp1dIRIltU38qcl2PMU+XLzBs1kk8BoBO83
2aF3lEBu4iSm4OjiOWmQDLie4DgMrBoquWQLWqrMwSSoouMgGtpDIsk4JV+d1TEEPhN5GaONkYgx
1ZLYW94ECMGWW/tVMHS+p3hIdWO7PYstrbdxIkmaLh8RK0d0EgQZzwJi9QJby2EgDXjLuR7xW2eq
gabXh1b7HV9POi8F6wrF9kIW5B7lVpGsXmt+MXxkNaTvh9UIT/wmp5C1/6I24XZ0VL2siLDED+w7
/kbpHRFq1xTKZc2toLYVFStsaroF7wiz4QEF70iruJ7+LOfTRVgpcI9TqPV7jxWHYTx7+wBfnVxa
i5gdN7xpTn7rvKoOsAMCseEYLQHUozBGk3gJiwDn+cdpFpfQC9MX2r5lCl9MA+wzZPbqI/MVcOTo
fUAsyAPc2kTcwneDk0dIm7K/MnYS+1Ifn2TOAL0ZAqNeAH6RfhES4Dg67pWn2TN9sunLlosA8Pli
2FNZd5L7NqHNCekfEZARBSJw44UFe37tXDMQXQPcYXJHT1hYlvZLJKDDP02vHXCAgqy4X+2Lg9qk
rW34vK5zurISO4gU+ZOndgl1YHA1AYpslqawG0KcXi2IPrz9Bn0TvUYqMnSq4f0decxjR4wBu4lU
ZwS+C1hk/K2gYHSK22VE3a+V4o1Vl8IQjm0XmnC2uaUqdjD2JBL+mLkcSwOrfK+P1kART7VAMEoB
Loe8tpYYkbKKuMfBe/ktdI2YxjBh0XpeKJtYyxPCGryDR3sk/LTc9pPxlMQriRjjUNJC1aaSsn9p
VNZC77aG9FBrx0hXfqEa/faoC2J8tjKIefNyYtFj9Lgvb+LwCBIjQbATl2WNEcPrq3CyiZx/pgZD
iRJYjaGWDG0emDkmjUGo/N9M+CboU34X47hbuJTadJPGGkFkmiswzkR/5lCzWqT5aCTVMh+8+7IS
w99GZSwEXKiy3s5nWOQJxeXK6wBQjZQxM0TPn+5lo/GWbeWaiDzjAv3SMwQg5eCTlRsDUSfwXYOG
J6Gsws51fnUdoJmd7IJg1e8G3x/jKtLG/XCvC0z414dahHytmAD5PFZRwpnEfblEvz2vQkZE8FtZ
CyWo7L3tPEGnoR+c/GQ0kfKHW/aLcgbqm7Xg0uvUND8jtwsPPUZ5SRY66KXEyWO79XvcHXdp6T9L
218RHfZdhvPfIKQSqQUdc02b/xUyLqFUxcx4kZY3gnSyKm5//3K6PpCANJ1E7h/Mn6HKzfh9Aamj
oDEJl2huFkhC+ilhBP7fVAg5sZd/0E0LG9LJziVjsvb2kQQqMSkDkjmZISX83+UpzdXsjHqhW7p9
xoVLjYa1HFTsZKQeaycbskX6JZBkb4yYSWaOq60TwU++UrxojGe+04/vEl0FlA8jk7nmAIzqteLz
G8krxT6Fmf5TawymUSb6VNrlXsXhoIhIXA8tUVEkR56ERr45Zxt0xH6zTf92w2plRKWI6We0pnbg
lluQ2HT4p5aiNUIRDKkjHrZOxNiUWaqW9/lAfUNvNmgyODIUIDqfoigr0EUlNiAbZnealwNXE2Wr
7wERGwe5sp3uJF/UKYmRQbcYi/UhQUUkqN/WaJzF2Lxc4Eqhc5c5iGA5V/2YctyiwroEToK2dpnq
mDcyTwhTbfPJWe5IvfAAEzecXpmIwpiGTr3Q+e3GHRuk1fiBZ9YoJeGNOXSugJ1dzFoKiqqZlSBO
ez4pexPNrXttOCeynROwoeCZ7wEo+e7fKIvZXbaIOTtfDiwBl1UxzA0IEkpnB5YpBF0zxSNpwJej
VxfaYj4RmNECA9zBsNpzA9ziGjz2ucJy7fG9TJrpw3Z38IrSHaztiStJ9InVGnd0n21AHWsvPrYS
2lm1+k3xPdzndIYHdj6+9Tq2/FFSd4rYXaktz6FVr/tNqqgSqeNWCLLp3LqKQBZn4tbvWyvpkkAj
CNnNomjzDelZWlrTkC5WXgArEXOZcdcB0Z9drPPFDaQ+sSdo6vjUViSqbmr11X9uRCJ+/TIhKd5M
LC+IMF+2RAiQIHuCDO0lvXs/HLpxLXXJCdpf8pgQ/E5rrI+nda/WS/5fCEdFytcoX29BCcJMdL0T
u0WZnoR9MmmevAYUUUqa3bNNisvyBVXgspcp2eoI3AR7wv1rzB5ywkIjFuPfljv/zGds9+mdKM0m
lhTHsIR8TrXjEnjljNBjeLZoRaCnBagceUlILdNO3hxTLO+R0xcvXWGHZMaZj10JlzQhqI3qnwnh
nytdrLn/A3iaNelyWzCR4mePfyyjZC9tWSRM/U6dWfQgKjNSNxsPa01ZAJPON3EWXtkuEYQVOI5C
9nt/av9fZ5EqechjKR83xGBrIjIaZ8TdZUOERi+cs7xLXCsbsSceaJPI/nYab1DEKwWegkSVZmZU
MOMbPM2aQV6qLnneu98JJMYnYCb6DXFV7QV3kv2ZLqXhU5ajnR4R2Mmicu36L74MqWLDIZVaTuev
APGQnyT0+AuYGXWm+0N+S5zKDv+uWtMUcSLXrM0e1+Db9sBPExbPc91ZW3MlQVRoL+J3YlkYietf
2BBr9pBRiJw0/sgn9miytTyMEl9RGcK6VUN9FVhHDu8xtOS1xjTQ5N+xmQ5bC1a7FL59aW1bjzdK
OoGvwOtwgW3kNIThpbCEMkmYu4QyzaoL3Tg8pF+ciLatR7sVVP5hMhH7o3rnn74A8YRszz6eLRnd
jvdlnl5DuA3ZCsQyZxS2RZWAHmAqjSKfGHamf8TrZN6Dg1fh+wd7L59JR5lWikVJBpbm1TURZ+Ms
gK4Oe2nAmk2eC580oW5lXxoY4tntasT1OzIm2FiFanx01hMXG6qntky6mM6mZe0trm3Ikpd2FYb6
vysdGd1knArR4g+0L2vEq+l7Xq0H5Ocmbw91or6nqOdMxuaELfE8/sj/n4IrhyY4JHcKPbv8/K3w
g5nBI4s9zomOW5XzKVtt0jQHW1yZgX4eXZrUT84ylMTUcHsu9NndLuL8ja1zrAZdd2+i303sjT+t
1fUva3ZJ2FQuB3TtXH2OwX++b+P/TLzCkCPvzwbbXAGrFZJAdKuW4dkBDBruTD8IB2ACgjNi6239
96xY0KQyWiEPbtAdqrCoG87884UxHBZq4A0jTPsQvFEp8vxR1TVTs+NTgipuMUqmJS9QxIyfLV/R
I2C31wwlEcuhmM9pWOp6VmfXg02Abqu7HsRpjw/dzK0S1F/Aa5bfoeQ/Rq+zQw09smUo9NrTlMhP
tyVod4Ba2MqMI11rbSy3Oe7gXF/xURCmB8MYrlni+50OmhoPQI4n0PdncrUYYDoCO/aF5cSd6FPn
z2jQX9kxmsaAzZRS5OeSAhSnn3ExAtE/rF653nqSjY/8XVw6VThbSkNP23B13VRFuFoXWdfN0rpu
LMG48AMmFVgWJxyl5S9iydIXmzoHWgJi0oWcil6/pwgnJ4N1RPCYBzSYOXwhYodwWMXCIlnWP2r7
NcA9dcy6zk7W+BKQONmpHi0zRvaqGj1oZTyq0QDboj9nF1f8dFMNH3bfJhYalSsmT9FV/j2jjth0
1LcFrKMAo/lQmWLYh1AFoIMnFy2FrsI0CZ4RKO7Fs7RhM0WmdLoj/WnPmXEk0vfofMEzdGg7FRHb
oRWKFsLxBFFa5uORqEb/0TDwZlD6UDb5ZsIjAYF2YYcHBpcExGU/JHD7K53s9z4CxXZ10zeR6nhe
IAfGuxPSBy8qb4f3M3ZuU3WyA3CtYrisKQOST7scuPZCsA4oyuHOPJGNnGGyukODKvNWkNZw3oZb
AZdatNOj2Qun/uAdbdmawxO0nRAEP7AzuuVD8HY6XCIXX7eOwoa/26zqCKHfjmAQHP73CdxSIodu
+16U3F6Ck7vpQreDn7kydKN4/NEoML/XozAvlKbSJERGkXIc0A7NxRQ9lVlDdtUxtGIp5C38GFDm
6+ep+DR4Jumhbpkv0h5t/EWFKDrksmrJVYlRYUl9ljWU5YoZx4JWEMnQwobE/LgBnHeyMiXtd/ko
Mj0+DqB+xm0ZvJEV0xzs5A2QOGsWwvxV9fTMD0DJbQWsEBw+F2l+9e/B0lo9h2ULiXQNg51LvpWV
sd0m7lu/P0hOvUgtISMZOZB5ogVlqZxuYNm3CuuXMbuOTLUasRNAIFPdbsKZWQXdnU/ibWEUreLg
o8/ht0bwYcD5YPoopLVFUdaeNSbHLsiv0BnbmrHc05S6lAFLyRWlGTqYfpwZjQk7jylQQK/HVVTB
LxZFnOqJ0giMUqh5TjVv57R+oUC7k6Ls9FFXqJQUyTuMRVH/w0dzBwKi2fHHvqMAltwPce0zjab5
+tMEFC0nif9IeQ9RJY6NGKLYkrU18t2p7LP+FpPyBm/L/VtniIth5eXze0rPeGubFiQmzNT0UhOP
XrEkKtUNRUPdCJYR3a8P4Ei/2sYXhwliSrJN7ub1QGhX9nXE9E96i0v3zB3jR9hJHGtbulnxy4zE
pSHkqZtoD/Fli+74w3nXPwOHFh+rnMDtFT39zzLWHfBLSA9dypeX//Jwroov5UJS/+F6HbsOTEyE
kL7ReV8WMUBmMKNnXQ7ya9ynJXMb38wT37KwvPrgSrrgxu/ORfsHZvUBlmanWKSlsmkgvPMOURK8
bg8YMcBSLFq3db1f+Vzftzh4ETXQwgKIznu3j9KwsVQFGS5PapGI+C8mDN50zpid4Co5fWsRhZyE
6H6Eg3LtsZJAEw+ZIo2y8CEJA6MkEyaHQNeKzg2yXpJ0hy/2Ywe6IVXR8hVh1kYlB5f+Rlhe6K4L
Tk7uDhFTgBCKH7ePaoFJiHgChNM71F8fV7nBq+opZwyCNy5huZr28whmEAQy5wEYRZnCYAhm+feO
gCfBo1V5KzR1ZQHEQvMxikO0MMtjwl9kCO1DKY4vqFSDTkzlBV8gsNIUXsHc0M7SkDcfCN20TPFe
MoMBabvrybtRY7K/SmZqFDjzwX2D/TH/EyoVp2qKYGM7dFNi2JoYWsApGDDexZjTwlrvitVwr7v/
QQljuTfwd49on6ngD0sSLdP33Yt6BCcW2xx60dN1TOpfP8yPdoP6GCDa1bZ+qTTNmoeytpTNN/2C
5rhFh+6Vzqnxs2etv/SBUrMrrMdecLIzU0WjKKQSWeHhHftyyqNt9w9uhVEZ2eWwuM1ZX59Rp4QL
/Y7PgTP2UWySqJpW4VuYFlmzR2w9pYhEnjSdBNywGB1Ix9qDkEg/z+DMxhuKhx2umC0EjjnfoJ/A
UNWd3zc8dPfddhSh+D/psNzZkaGtq+Zn83Hy6U4nWQPioEmX91NiHzF9NkjSripu/7Bek+wyj9dU
66U/N2/Q3KVME3X6dR+Mx0w6gzuwf8wAuqHcT1BvrjR+EmvPCmp9pLrQFbxCK/UQguzFW7d3nyVv
pFuqEK1G9KMnEvNJaOxKw/5ekCAxoPkFvdsp7CUsfDM+n+jLfQHaIuzF8AxLQNRSopKkwS613/NI
oXRJfP1QHLFkFOfSa+/5LjsS9/BOyMNxHas1lvkPzgAzaiVq2yVsmK8dHLhF+aluklZQNbm54V6p
hiuMlrqKNq0h0j+AiwaIa2MZ7O3ya7zzECRME7AJVVNCuEu3fCW3CL2uSCOq2aE2cpFEkNumXqhV
31YLVwfNceb9BhTxR/TryIytgUZ+lJn4+joig8XPPnnzauYjuPcaGEHp2vAgvmWjKAScIdWpR4Jv
jO+kn1LWYoOJ7jXQoMSSpGkYO1d7ALs1bHUiunZgHprgAO8H+ddhhuDbzr/vJ1WxCl1J5wKNHspC
39nKajmJZdgikrBsukt8j32llV7st/p4rl5chBNu060FJWkwUTvd0DNH3j05LW6tOotjWwDN2wz3
IQxdBnqRSePxAO1cToQTIQq/vnRUVGfhpQa0cdFrEeyJglijri1V16x8omEpxNy9aymR/s+sRMR+
y0ev0UnUWh1nqWP9hrTSJn15rhtpzc5kC/DCZdbDss0GKZG71DzGK9XJce2MqpcVHQwT7V3BJBH3
TXQx+kFvD9HyvHpvF9mLnwRWPnzAyYe57ovH18o19A05YxzPltSQT0YJtXltjsP7NqKRMbnO+OMw
WOhDJWtgpk7dfBnwawKFestpbFiZ4JmvHjIjeIjxfiVrWgtXIDTEVBSs33sHvpxPi8Yaw0qGArzE
bUMtjDHnh/azsPqySG8/F1CNpuSlqxAnW4cQW4p0tTtED2zDCdpzaOUc5HNS3SMEv5cVAzdlsvPD
LR+ySqobGpRNRptabl1Szy6+w3uOdNwlmp3xaIQ1cmizU1/xaDTHLiXvT+YvN+AomS31mqiKhtXJ
i+LvoQfz8KNpuw0D8Bq11Yr17z0zU+PxNs3/yEAemSJJGBkD4h7CS3J+1eLF4SeevXKrku9V/U/R
mgLrgq3LfxPbFXqkhB6moyNRVEl3uebL5r/C++kD2y1niLK7EMazXYyf8gNGSxeYgZ3cdDt6V4Hs
OvCUDF54e2BiWGsAHmGRQadQaeWQSjbsYzlaG6XzE3KL/A2wHKGj0iZCKmF2PnhJF+lIkm8mKPOh
EGm+VJTIlL0oqhpiHntGVVifWdjKh0zxNDJgrwQfAEMf9fkMRdxAPvF0z+v8mz1jKNWsfRsSr8Z3
cXXRJdAGNWdQaUviGiwdJ5Go9wzo4/MF6HqW3pz4grkYhibR8KTLJRTuviCctpjsH/Fpk58/2rwi
ltEc9k5ruvxjepkN5kKCnzACMMxZX6UKALwd3esUCKJxK/xFVyN77wRtnO0ESO73MHT5VUVlp8RP
s98NzakuiFcZzcfUEo/St/Z80zSxPIezhu/WO5K51FIVDQBiyuodd6sTIUW1Q++NZ4g4UHwtZyar
9GQOSm4LpE4SUGXvwbR85G8raJynETq+QcPu9kAxm6KSz7a4UVMd1TGe+tEzkR+6NYs7A/kCqgkd
M1RH9x8TwmyGjbKcP/JY/owrGJRsvQ2i6Ht/9oJidwghHbLMyzNOB7l+YQG0UGPk1b8PgFlYz/Te
zNIAJb5yzFSFNMdGGLyKh35qWRG4Br0PE8QEw3+SDcboXBmDOq3uB3zAwoFJDVMB9I1uap7/Ztr0
9EQJLhqoSFCl+l5XyDv0HbTN5/RLBNtQl07KpGga598NHoSq/SiI5C/2Co1xWNjxdf0EvBHGKWqq
Rt+n1Dulx1NSojwF5T8R7kzbsDbNq3NZ9iw99wLo3jr+y9aUcC01pYPogYRhfycfiE4j/Cf5FmLH
tLLaDdsPX6n5I56uhydVte5zPOEmgSrf2R3vCovehAAZSODRciEeEMGQBTg29nuqmIdnpmehTsrO
oU7tcF8vKfyKcpfzcmOwH1WVEVNMHEezysvwaIfFoi07M86OVGXjlLTZ7bCycyaGJ9nMbMOR631Q
2Ny0HvACchzgdpg4F/0zp5PvjaosCi58FMH/nSWnePvrtsHw4XY8WURcYCqvnrkMxmr9ImkcJ9zz
aT7kU4ptbRwOpWWgkVOcBJaQ7vY5To5+GT5unXxIWLUUXSm53KOTNNB23r0oChhY1hLdKMRCFFl/
QjBVvcDmMzxr0TK0b+nDCycQzcidHtLgiZ1RlQP/EYEDYIY0n15PWmNs43CbwpvxWgKXE7duldPR
EiLqTAIWw8WdTG7jpgixki5ZtidfvZJMNmKSd4nlX5lP5PWoKjePM0ILQwGTEzb2NPsuEso0inTO
B2b7CRbcJvBYJb7RwIIWk3BJNInpqShAIPfxOMIZhnUPt+2uvSfUl1tXc6G1T3yIIppb6jb/h/IV
16nUSfH3Kqk43kog+WQ1gJXuUsuNLM4YAk3G1DVX60uzQYCJsIpKDZdlHO/CPBqfsMNDzbPRktY+
OIFpPDadhi9HhguYHK8Yzp2cqJxEY9GZd50Aja6uYf6fOlsUq4fMvhwEtnI7UFfqta7Gnjb3kKI/
lvsMZTd5bS/J3nKctEagd/JQAL+alpiI4yBBSwuMeQq6FP5c4EnkPvuDhl6bGK4Der7m6BmdUWCf
HWjRX5sypFosNLLEsUCvr56ReI2awzKh/oR8ZnGtPHZpO0vRRUN4n0+uxB+6MbYsJOrB+NeDkfvq
WFk3z9G2FFpi1Tib5G9OmDQF8NsJNkuk9hRsPVNKojtNwcYhj6a6PzQax5YI1T6+0DIRV5h2aiLa
WDHgoUmLBX8esdSFdt+VIMSlyE3HrjmCeVNCv4plM1pMUUjpJnzNxsXl/Fw7cxETck9vKtKDinui
p16WLWbVl0KrHLIiYTo993uiJNXs3nff+k6xKPTyInPr6ud+OgUVkc6A8O2kYljMpezf7MKcg9EA
ARZfJ8UQ+JeMGNDOVuD/fgmdwjPuXuz24H/rlc0ebG8wpstEDP0Lq0x3XuKlqyo6fGW1XBWr24yP
zH8w/SQkWV9bBlWoQxCVUsgu54gUdWICkA+9FpDbb//SRXz0XG1c7fDzc9kAckhjKd244UwdQWX/
sCaLLHE4wvAxsTAwpBbTL+AaNp8qv2lZEMN3Zl0mvL9ihUsJuLJ+q0Y2Xv+rCx7a3q7RuNrn2DuV
kg1O1QCC1OIpgJC1UGapezEEM3Dc2EAOgCXbWwplsMgfAuLoCDD+ARF/nAZJCvGzR4AC0r9/2MKL
zQ+ffkGPQ9dy5AntFZAEXD+nokqKoWxLNGcenr7Tv4kUBML9dQzDYKRd9SAg30u9m7uQ07vyFt4M
sbrM6M2TUBWmRuN4SYcgXSp+TfYcha+rSDLGolqYHAsts/1ngZfiljH8MCaaH++N65o1UtSxKt2Y
0gE6/KUEHqstGiZNrPSOHLH8FoUzTAMjBOAQ1cMijohjgI2WCaG2sXhALVJkHktBxZ5QEnwXCSnM
UqsZsFMvVBXQg/Gh8qPCQAoTW4ezVZ9MVsEH2suV0FeiRTRzqSAN7vLKI4I3ip5O/na9CnJZG6Tw
jZDaHSgCjl/JSrVX0IMLhmkGJ+aX640I76lIS3c+suUsMPcynfGql/J7E6u99b6hCZ8166NzSdHn
46H8Xe2LVD2nPzFRQU2htAajGyxIAgcGoS3eyyMkObHp0K1hNKp7/RocFfpJ8QjrDLE0n3sqB9zw
khZP8qMXfQbzogreHHX+UuXWZJQ+Dffp4CkHxD0O8VOPn50HeoRtna31XRoKWkAquX5TXuNQ7/cd
uhsRYCj36bG5lGQkqzlT2+aBNTqkPADW2fqtuIaLIPyMv3PyHm45aPEe0je7/x1u8NukLIPMjxFg
tXme7Zju+v9zxi7rcnrD/uHNUeaOp0qQL3prNlHtXWxXj3wdvQXmS9pbHuZMxvJ0d9T8CGyz9vn5
1moaIDLcgGDUQBGlvm/6lVs7j65oWpRRfSbzaomx0wuN1dmXn9X7Wuf4BNX0zOt85QK/fd1ul0OW
Y3VpCMwr1irbRa9nV78GnUwD3IZvgYtbvAyCyAUD4MD4FalG9d6sZrEM6D76F2VHPmrSLgUeIGCU
KxUY8pfKdAUF1jo2gQIHb9m/7Ey9fhKwCpCsjIPu4dQJT7t4WJNTmORDdWlQv5RmNFRBgEy5r75Z
cAaCnSWnQmuulh+S4ksk+L3cYgqJsV0qR8skoAkN/5VJ9n6XCePS6/3bWF8VRhUkcQRrVHvbDQ+y
akImFoNWzDawbtp3c3Za+j4EZMkePe/ZoY5eL4ut7f178LILbAi+dlhPlvjvTYW9mLuAWdjIMtNx
nKognB0iFfM/oVNQjVSQaOoWVnAMXKRKY+VzPYUhXElyC/vjbCeEnoCgK3HSj5zn/PJ3vRvcQ6Iw
Y3EyI+dUHkKPyG1Qxud+MDA/LuvgIV4OUVo/cZfLU6TRGzkzy8ylGb/YDzGR+QOtuzer55DBW9Cy
Zr5vSKx4W5dxcvCDa/MEz43o8wx5c9cO9g7hT8SPPnPJ+Pdi8NZP8tkV/lueCfGP/uVVcqdTIbI6
XzCN2hhHhOoFN3/pqgdpngCKWcZ2/O0Sq5j18eB2FIPfECV6z9i9CeO2O/5/ac3iXJ/kVSy01jcp
82gLO4IiWzWYXpoL+pF8nr7uNM95WUjXisrvX4pcF0gCipbelfaG1bEC9KnOz3td87FxN3yW78vL
Szho0RKpcu++1BXt9O0DRCIAO1+7/QAlPbRG80c6hhRJgfAVwcUg1gOwXg8bbYnkG0MRsj/YMfq6
MwLPts+zpFQw2BlDtm47G2Q5hj6aJjO/3h7jAW1S4COpqmwehB5H4hCFVphAaYT/elmh9OuV819c
WqBut6ZKUtBGhCWsUDiRzjvhXwdpCJWnkRk49ewBl7ZWftaYZZKBfjZj8yFYrrG/Pn5dSJGd+N7I
r/+3DUhg6bfvXkE7aObjJ1FFVbD6p2/gotD6qFWW1Ts6QQ3nmtPP0Lb855AjzjKsJdi+QXRDyYVK
nL95Y5bMIcLicLcGIfpTuzmNb2CgDy0SjfJbu6irvOTkcO/A6oyzNmk7K3nTz9SGqKoSJ4EQHoa5
Cj4FJ/mlJez55SMhhrLO1i0KDJ4NOwK1MNoSOH+mCu5sX1nHf0u4sJ2VG3GR/lDfMOTB4M9ETU6J
7kOXBbJ9lJY/aGA490+XFIQ+FjMeShpuzcNdmnUlG5bN1wre0gORdyNIOVwkwL/b1ORzFSPPHLJo
s+XRugBXkL85Z/a0wtQ3ciiDv0wkVTO1WPBl+hdFblSQ8uFG0paNLmPYghBDbFODg1KvcdWL2aqB
StS6nkxhP270scc0Cuapsrtlj3J4zMAh90z8GIkUK+wtMx2DwUgYUSzD0VoXnk4XdKYRa96B1jJc
8BxXrLmO9I+FW9E0bUr4AVs0Zc++F60smhtrM7Znwh+zEP8KrtQpJOy53jYMCwVnB8jrwve4fU3r
gAo1dB95GTiN8L+BB+aEw37zoF4nA20PXwDGjZjUiACdC2g00T4pK7fPyHbsElceKWjmTbJRkmNE
E3fhl1Iz55xF/wGtwQ9KNgrPDv1fp+yPwx+cgvhYGkPrUfcixHyKDQl5OeJg4H98jUv8EQOL5kkR
ieOH0qVm9C29g2v1MkEH/YMXLAsjWXTMHBk1u+yOfY1i7cPbwqiGmrEyXBSTqdGH/E9maMsemH83
UBsJhzAMwxoYaANsRPb3eQk3eDXI1z6QJB6wmugr1nQ2IEhG49pBCeJHPuWlicln287TK/rTIXIk
XNiPz5mAVTnMnr0kSv1uzVvPWTmxCnUztXxU/O3lS/AKrPSy/O4gX3tXZQRFjrn2qb2dxFKBwU7K
Bb4VXLXLrImQguAaLfpKzkGOcmWtGTUs9tfmd8DOsUmUTjNc9T/eAFrJvm5oTYbWHGugG4TR3mgd
F0Wo3Y+RBOALAez5n9GAE2o+SlSge84GH0JlVphggeqzocxQ1YWLYMraPlgDPqHoUABH0obo02V1
gwfQcd+cz2Ril8TNxsPCdVF0GvrFFPRZSsZiX0cmSPFj42sKwXAhPA/K6qnPeFM1+QAzF5ubxQlN
KGDN2ohKkosnzpeHuN2Kt5tmQCbwIYqtziM1JAvyUDvtHvZ824l5SsaZRx8dp3UIoGdOcjbTq3OM
zJUJuAP7yGdKAJlLENoDa4eDP/7Jzghq+1BOG5jdNIW2ZH4SULMI5bBK2Qa/KUiUfhh0ZnSDv/EG
a3NpQAJjz7Xs9YPpNbx8T8uoEEcbI0uUqSiM36TCInBkaMxXwOMC7V4xTxh0wgSSbF8BgQE0qhQl
vKVaEtn2dFGTmV9/yxrIzUK9e4DA4rS5SW65h7jHJVvSqNSTTm5opmNUszPz805vedMbRJIZcJNg
NsCeXVPQizRpkq2A8ozy/RsQKHlmruOcxdbruxsrvDhHOg6HombqMaUavdqidFMgflRtv0DD43Zh
jsRk6Lfx2V9BjCHeqmWypeCJs1dTZVUXsGBhfHm+BcnFmflSYOW8C1JF9ftODw+tzp8cQFkCCF5H
31vLx/w2JZ4fHzlXUIP9Jgu9vrdc9X1WG3ppAZP0EU1dWXeToRDCSNyS1Zj/i05tujcB1EpDrdIC
o+5cXJdAb6YJFai4U2bA/GUQ6Ioj/gFczii8tBPhG4stqnaLq4pWcrUNqOM0eTEn6kz/oY/ZJTuC
BO4u7PmTuFgyuEntVwgLB/qzglKhGDw3s9niBXZKwTiHCV0c/Nd0fiB/ovIERj/rTWMKISBSQGIy
/Tdz8oE64z1Uwi9HbNsJl5eKr+OuE8xVyibI8q35nobxqLUdRLDGfq3B+d3oboRa5TFb/rD6Lnru
yXiH5I6ExQoyxaXxgRR32TqnI8UWGwNQg294vYdrwCsKLS/DO9R9rIC9YH/Cr+pe7hQeEvOUI5/x
t5zaOHKZIJe0KBTTEDyHxzkKIV4Um/LqlAnlRwe90NlQnxLgo2hkDsWwLk/q0ClS0G4NaBJrbT2V
iVcZmPIfB5eQBcrgg3+Bgt3wNMk8JcNFv3bEDs4KDO0ftYuS+lpFtSyGwYkp8oA7wMI+KOCeIrd4
FwrZSPuVMlt7kQsTmTIuGJgtytYzaJocSKJRvt1hhfLsUv7hLDWj+EJk8whEadFo6Ghee/3RITul
Jdg88565OmUdnklmJQknlwoSjlc+ICGLJ5udyXvWgX63zPpY6q4WiUlQ70tiaLLokxggPc5aRmsE
vzu9upYWY51ZT5bAf8sP43Mjq0gpY7X6gDDig19AxjOw8uQutDoYW500gT+32ZUuHYiNNfIKl+qM
6G1ilIbBfa+2djuyqlevswkgwMAg2HTgFAHTQ5viQQ7lM17lkiksdmHwdlLkj7QWT1th2rcyZlCw
70qFyV3FTsoHJQdShYyYtNKYlsIS8AXS13FGnoeJoW0A2WXsFj2kxGl0X1sPOdUfsRkAsSxtYY2g
KcFk7NB7aF1sKlZQWjmc7/KLNmixwHqOPsTHlxZX4ULkPvuULyAurNREboShGphFK7H/gedQG+FO
DSd2/na9OEfSTXX6wJefzXdQhisM0YJZKPxqw5JYQbxvo9HUZ9funTG+eUdn8gvs1PHLqehy7bBC
v5dmbxJx+r9lSPY8krcIiDqEicjdlMepcoRsnWMlMfbf46VANwWFqVRMFtdacXXarjo4G1mwoGI2
htVjewMucj7pg60PNvdHnN+3Jpjsy5gU2bDBqxAUQL2L3rYocFohczWiPCpY28zWVe+Ioq+iyspq
Uxv7/fwJYCk40E4YqMWnqWOf6JYboRYL0jQQc+L5DbQWSb6wGbjIv6Dle5yUPOLvSSQkbeBg7goM
VmyW63/SOYhvq/XzExKvYhJfkOwjl2j9QcluRSxcXrHL16cSNTjp1d0EDptlHY66pO0LV6izI7ke
YPqHveG4xCg0x4Fs1jeIsJ7ggjvWFsrbacuDdzor/DTvDsPcEUszUVRvp8j/uW/bMxv5x41jmlJI
wBwkwACeizNc3ZyrKaT1xjbXrCMbn2RVHbxWd2h9iLydYfswHfi074ar2hUKdthjoXJazu8bn509
4hH8SvNUh+lDm4cW6UM1bjJ1N3vu93goxTHQoGxKPx9aCUYc/vJnZMZ6Ylk6SrrwV1qAMvdU5NYO
w9hWvdgS3PCMM8dbnWsEkNkuPsEhoy8faF8RRou71VJI6P+vpY7cZWPSM8PZIoOh/yoqF/FlA5OR
rFEXDTujly8aKGM6YTgVqYtgIZs+HC3mpBRIOTXQL9ME7lWfHVHsLVGj+Q1Bpx5ooKW1/SlCYGiv
gXaYKM52InpNuX4z7XBehpKftiRGDqS+pM3fPWfjiNbb7fbxo8mD0Jmu4Vh/c6OtxTQ89wTrQOSg
iPSdG1d+wqwJIMrLPWypfCfBzAHR04a3IDyKc11FGVSvgM2DD+o3wMpE/zTPG0SygjCXrnQIepAm
MeTL8j8WizgQrXaMqw6afLLqK14jFuhYn7V1N536A5UY7I1DhSJN7pTOhnQ2FiCUx9EK+orTGWop
/3ADQqk6MzGg7fy0jqrNPczTZ1/QInKOuT/dKimBJdDPmXAwamebrWel1w9fx2AtcBA4cMRwyd7I
zCleAMYGv3nk+dbWMYrNn2f94+GzoBYonRFSkzAvU6n1NPVdz1CubypcJ6uD3WadUbFC3AQtU2dL
v0lXk0gzkLbblmO/HbHNLWDsEwBWmEd3FtdLpsDppo807RN4wSFAyZPkWmwKECxUsyJMDKr9uYan
PsjlNnVXTTKdUNfkRo2xRyXjsKzbDPX+UgX+NRHoI+VjHq9jk+XgRME4vteIeogZfjkx/osul9H1
QqOJ3VlEf9DIqhPaktvDQB1g5bchB1PDGN0bSaPvHiyuPt+Te1v6d+NrIi7AhUnwBoO0xJyj8NSV
Rala3n0T2UPxVN5XNTNz5EOzl/roa2UdOLy6hGhDxIMgdB1o3auB0vjRtdYXKVJc6FAq+jDj5jhk
8xuNIAdHCzNokWpDxzLHm011j8G3ISpA70VTJZFalVM5O+VOZK9h09aOyaj4N1lbaV09hqvdXSIM
SMdUHS1u5o/Gp0PLsYQ/F85STncKyDNBDfa21pP4jdd0Qh7lmmHlkzbW9NtAeg4RRvY+kVnN2WnE
OK1gcIcDzu+C2MdTKqeHmyX+F948jdEXnfiWX59VkIia7dO/fFEVTLjGnPaCbXnUPiUsEjIE5D5q
k/Q5Kgo8ZOk+bG2JGLmhTZsPZhfkd6fR4zGNznlbeuDRn8joMBjh/+RtKZ/K3LOEtHGc7BAAt5uL
T2Bd81mfqC1Dn6RaLmRphDT9HKgVaAj5XbsgddKzVnoq05+dFPcJrxhmxvpu3+4KICgHxWLfLFJB
357EFkEh/P9+8M1VIy3lz7yyvwvPy+gds2zXyXXHzZB6eWK5fI9tbP8gMea7ZkiYgDCIQWlK5x3H
gSFCgAUJtsG2ccQcdt0MezIRfZBXni7HSf/9OG0uQ+zKZTSB90kY3olvfCQvPaW01HUTIF0dKLNx
dRTVGCEOlfzrj9ToOwO6/KreDxYgtnd7rZeO3skO5VmbVKqOojTXeca7k7llcYmzNro6VGPqTuR6
ld4Y+2K6Nvbeck6JEA4QyAzSeWrVfnZnXfL3mHg11nQqZ3nvCpaFXlQN+rOQg8Gvgfhh3dZzmRwh
6FsPhq27i9QA5nB7oldxANUvbSO/z8+0tLGD0ll/PJKHymstxtlc+vcj2uFKJ9YY8cGp19fhrXgC
btpkO+tLxyMD2COfPVnFnS3OprgJHedraYaUiB0ZVlrQuYSFoBwlzjAm8SPpBGbQNgHtGSIdP9Ej
aR/v/5yYQlgfTvaaZN8wAK+9y86drGbs1VRbwSW2KzFNxXGk2kArm5oi5K7QHzUVZf82Svg1kd4i
4JE6Zrw4SkijdjFV2IPSjjWn5naZv6iCOPNaAsspbBHjFGfscsvq2azVRTJ7/ylvg64tBmEVJqoa
HMmTcMD7xEYcoyafMkgbdN9tJzqnSoPsD985yQspgZd0A7Lkq9Pao8nPVpMuryImB92aAhsNdBrh
LlqZVtBvKHSK5WGq04qqwi9GeGWxqIdqx39+6skcNf8JsPEgtQiKGK8IDr3udJd/yRcX/GFBaaV6
b2hySw0V5We6i0sabhqs1emOHfD9Bk942FWOE4KkF+mFQi3ypDu03Xa+Ahml1367mQuKbjbP1rsl
eRxNKUTzD41Ez4iYCIW5zflMya2jyPpK+1xWA5LWXadrXekGzLYyrThlYXzc8opwPI6QmPSRIfBv
0KNSLjKR0mFzNjHXUdLOFEyRoQsjZnBuUKgn5FQYB9D1QQkLQNC1qnx/30VSPpvt11YBUpF+4T3Y
H60FninxGbPaXXHT6OU7hZ+0xprvtLiNw09wax7Ad/+C35HeZdAKXogjeFrOS2CQ8/+T4c2YUKbj
1tKkw8/c4jAUI23rTpVc37Ov3D0aBvQ/Xp66NMmEuYhDo1+xT83Lyett7HslcAl9kRMlKm+6wlh3
4pvsMT/M0UEDh7XdTEhahBrpzYcGNsGYFA8vpoXaFKmE623rM8PPJgIxm2rraxFTEeq7pp1ubNAL
CfHcDpqdxdtFZCM3Pamoeo/UFtaH9kWOVN35v79R3SyfD27SNvFba1CJRDTguC25Pa698fHLUAYT
XhAWnRTGrHjEqwff7nJOxfQ2Kw6WfbAI6J2+yvC8gAJNveGu21JOav1lkCIlmaGv5yA+cCJxRVzQ
ISklE7DhtJBup2c+7hfMpSkiZgAKJicSgWNR1g6gCFYlJK4vPqHk2Op5BuCblq6ytmfImTgt8qLt
42UUWDi0tYYwzbqGCkBlNbhay1G2kXL+PyMHg5aBecRYNReDJDQX3Fosr1YM67JJLfnQFaS9aM+0
ACf0/tIOgMoP6FZjAIg1ElmYp8yu8bHsLXFlNwfJn7Kx68jcxdoZzLgEWU/7fZAPOqolSIXiRhHI
axerHkEQQkMmezBSdH80QItKqKikK1rLq2wYiR+V2GfTw3jkVza/2KOLxPFZmN0X+jGIL43DVg77
rs/OlQl2qDAAPlbVXzLlxq+Psgqa4UqcQ5qxdQX2EYhTAucRDDCynRN69HDql7WSq/35ZqCLlZK8
s53znq8f5GztM6bR/s65RG5QwpgpqhKq4FLZ81t2aq/OlSCmHlK+P17p0vwHPvRDNEZHFr6DCEsB
wn/ee0e9K1PYcj79iTNRLsrXkrYgEor9aamGi/HFkAY9dJAV4Ge/Ue14cTYzCa4+h9NiDx62knCi
UINxNLU7Fkt8kVRucIpfGC5soc9mTaD1ojYh1Mj5LLyimhO8bckz4ztmEA70yXqz+JlYR/faCHZw
0urzWPiDbCSd489u4N9EhcljyF7JI+xd4lEWNXyxxqSf1Nh6vJJ9rk3N0V8XNsd2VMlTNBfbUBEl
RzFkGuvtPeFuWbEf2s3jfsOADhV2gKUxTvDCyYql4rS9UtnutH2nvrBHmYlWcrC+5WGkxRH1LlpB
AAOl0iRIPdUxFawMIr6N1KLxThmpiJVc596NCowOGGufWFyMF/iGvSaF956AcldZJ2IwoXaS5qf5
akM6YSi+qSJuZdvkAjIC3ncmomODrRh3O66QvRmlHMLZ7Oig9xZMkOedIFSFYZFFRZo3LIQGKU01
ajxJoRmR2OQEa1UGKtMOapvVJuQtK/3kX3n+sGTK9EdT2yZBCWGEHmmuVliid+AmF7rIcpz3s8bv
m+0IRKsLn4E2h72BLQSc6sM/iiozgJKbR9Rf8EkIaIf8v5Pt3gh8mhBN0NXy+Y4qSeT0ALMpJJUn
qZMv6JDnicSDcbNsUJU5Pe0mqe42A+RAgr3Csa/vEU/9sjwcE/wcSZt8sVWFfvOY4xaRWZGm5hat
A+oSw/5qXOEJTuQpQNeNSMgrA6mOCkkrR+FTApczv6hhCSi5fvLlGZQP6OBLSS3YtPCVkt6ChQCY
aZX4Kcgx5RS44ZICZ5QvLBuJw3/A0znzKCgyWzTYHFeO+l823k3+ZGhy/YxSuW338NzkSp5Gk0Ri
OHWCQ1AYS8A4AoDPcdLDN/rnAC6BKrX3O82by3CSnmzzKpcgpOR2JAJjFsAiTbPP4+Fdfmf5XQBM
fqsG3xi5RcuS7mbMUYOBHosy7hpFVqal+CXOj3KjADRn5arlbFcCAq+WaUkaX5arcQrR37LOKHAg
C/rUqtcmExmRHR5Qm9Li++Ca4TXUqeIPwYgE2XuHXq+a3Mi4GIOeJ22qHKZnSTmi0uqaubL6ixAb
U4UZdfJ8kCyGxeFnfsD/w4PI1zHppCLChbcLltgw+BiweCsuC9td5YWprmgKYT/UhCB+1lKdqw0x
HCv+PbFZG9Cv1bpBd2euCx+BpQGGvwCM0P1Tj+mbTlCj9jx+QSDC8UOKgUcwVoP4E/SBH6LqWzY0
F6lUN3b8foKIBTxanKxP9juicSC1sZ5EDlHHkB79rCw0JVoBLoT9SdqtC6PJLXpbNwpCkGrlAX5X
8xryTgNaifxDij7uWHd5XEdIBU1MM1gWpUQaJxIIswR0wtH6sVewSuyEJxRAK+sJw02OdRk4KjFb
kvTR8enUU9DzWGQIGeOq4FPs39YV4rve4UpMsVrdY4Y3tqVIDD7cxydTRfeweobXz5jbQ+DGGOlN
AHsqrGao/cFQNVUkRqdB3gPJgWqmg7rYN+6iOpE6oEiHF6yFV83zQ3WvpNeJkB1n60j5aHTnsCVX
oxGZYH/mSz69anoBek6jWSrytlAQqinDA3lCE9EzkJS9OjEQvPrd0U+5EDqTgAiYCFdIDygWvEQY
bmDGgXVAyVkmKZL57WwaCfwraSDuV06Dl71O3ClR2D0tLlFXpOUn4SA7M9KaY+jNOfhKNidMKBBz
fGlWulnx51L90OU31XnyAkeLOdoqZfuUnkpXEYCPz5BK8DYRYeNYlGgswLFm0spOXeTWvjvUBzT8
R7Gdza3utvX4pWTjJim8OuX9ppiDiZhzubDcss37AlaG/kv2EnnbjSo6TzWROqhsohTtzaxxp70R
MrO0w7i/he66yLPbaNqbxzDcbO0j9BKWaRX5GYD/wcpH+mRAM+KagxR9JmZSmdhEUloXURicJos+
SU87e7aXUqtFZYmiagflCPY4+GjIUM3BFoYN+38TTYmvWvHUd7ngmtMpG9uy9INo1smNsDn5/jri
49z0aZ2qsED89ZnCfdzhyOhnMIKthIwzZcSfU+ufBLJxOko9W5fEgx/zv7Pj51gkYmHqreHB43i+
79reCIifj5DeyMBe4lNm2ZyQeUbYZO0D9HnhuYGkmIT4hjMGPGdCRnOjbsUEXuuiZspbt7Wa4w9W
75YVZ0mk7/SXna9/d1Vnzb+sm+O4S/1JugEJFUoQuRRuW0VwHbYX5Pu6WM/YAVQ9+aiF+tVRRHQk
AvMViF7+r1cX2UW4UJqZMcorwrkpfDw9u8b0anl62yRDvqTDP8NGXCeoSglzbxmZxtmic0NDKw6g
rlBWA0U4N7syLMXM3zTZnGL4V0JNDm/H3QQwjpHND4HfA3JY7bC7Y2RTtQ1cbR00ebjZWj2qP50F
Fw7G6b/Fkuh+DVdjMKFzP93Sba7ctyHaRWrE/0US2FC+LbdAFJU4tzLZ+B4QhEqEwe1og6C2EFCb
E9TsPzLpJ+mK3uCJVS+SEheHfvL+/EJq1f8KjSUbqWoIDnzKshtlZyWfCGdrBJlm09cD5q2gYiRs
IqiexxtsvsgxozL1q2Ffws/ByaMMWXtFUbdXyBSjhOpSO2g3KoS8Tr3otLzWqt40V6xYzbGoRfVl
JniyOX/8Bb7eSvg2MDVSeNWfXuH4ZU7V1awiE820tZS9LqEqIki/wZnhRZvB3TX0KH6WPmqQpCqd
PbCo4Bp9/KQwsAc+MbOxJW8XtuYTqrKmMJ568taPY2QQVx03IKr44ffGaw3wY+g+KeVInSdjW5cH
t2T184d1t8OY2qfwn1KPDxAktqpZa6acidqhM6WOL40hrjLsmJ6jSgWUMCE8b2hFQqWXUZUTMaoD
cv82mI/8gcQ13i+gUyXZtqJIJZrlcfKCJIBrzzgtW7etzqcmkoCLafrQvZ7aBy1rjNWfjtPuovMM
alm+Y/OvvPy3y3QCb9LzPMnstk5PjFX8Yhgowg+PLoAjm+5I251esRphG3FTqrgJhI9XFHMZQkls
x54xvbqWvHVTggvJfCPCbYOLCP/bcLRI3r05L8lSThEjIDtQ1ZcVnnf9fB6xiBOOR6LOpYWb+ShE
oqrNHNy0CYqHe8+6JptAqoc70zuh7TBqCdJIlUxhuL2mzo6SkOmjop5JiZbyzbhD2vHTXJkK0MQO
ha7lRvbND7fZDFV3Y6LN2DNXUA/AQJpBWtaZG0R4mpt84pKxx8Z0UJqFbFv0lSCRPX+MADCqCcVk
UNr7FAVWM/A9pn3vON33l+M1rrTPrWX8DK7yfwVZtqWSi+6TTOsuhQMX5O6Or4lCVDeExBrUSZpw
qIJnI8zOced7/tqH2sPOcpCGaxLEdIzkmy/vTzVTbHHJL3gQaG2j97cdM9QTMXo5JJoNxiAfPpl0
lfAdrXKr2q4uzjb/nHC3S7UhAvGRtt+315T2K9NU2yDa4aLEFUbAux6UJTzDddCYKqxBnFjJrOGx
YCA89ApSrb+umGEYog826CxN3d1guWcriE/c436vuOpuKY5RR2/ablDpNAoXZ4WwkcjWLePgH/+I
Hw6ojMJJzv2/TffzRVpU4fFqrdBRrJ+k+qjN4lEE8hoAVqEhfnJgjjs+sY/yuLxwo0jUCxen0Tzw
5VXC6krTrNQIF9VBTGDGI53KqRtekwb/4576ZggK6sKwOIt44KMcB5JlUUS7lvjz6t93o0hpJaTq
ADSgfKZdr8Jxe9P2UF/P17rsqZEs510Dnmfhm8pp/WZscHhVF+7tFTj0UuQg0CD2uoNWJgNvtjuC
BhZngH6hL5sB2+aec2uGoCzT0jhdqOrjZn5mI+LIjTurpC63iRCX5QN2GRm/dryV0/tQge5hq9ey
wMGBAo59jos5pZB0SJbYzF2P4nK/gDoDbRjJzMZUEtgqSbDdMP2+JH+VQ9LDjkhEXCrDbLRP6+jY
VSRwOlgfq6Tqpyag1/uWcjiwKjM66SHPT5c7yTKR/M0QQKkw+l6qiFZwP8knSrCSDmlSX2w187sV
oU3KPqeOEsumQ9qtJGR6RT2t5Ah3XogEkZ/6IvWwm76vAotTy3TF+phY0Q6TeR5aDRTlye3PO8aZ
bjt9BycL6MiO/giA3gSqOdMBAVMAhjBFif8OcqyyUH9GgTykH8tDyOO68RlSZWqiPyCe4iqoihor
A6JW/hbVc8U1bMbAmVdVGqkvZ3pYYm8mOYH+TQRm96DLQr5d0evHpgtF+E88k9H53i+VnpnBICXA
yJ7ItOrlBHwvxBUXAfS3u2ilNSrNQG2sXSTwarb36u0YE6Jx2q6fABZttBdAL15Vzs6QxTsRSYSt
W15deiZmeQpOEw8LbgMtpE6IKe6BM1tWz7qMWz+9FzfJqdHtPQteNrTCzjAJZ81nutWnRXHZsRxd
8D/FCR2LZj0uXm823iPVfnhlX2Ug/D7Am4y6xmX94/vg3o4beczajS8KEoAHL/ARalSWqTC7R1Xe
YIvOBrT4oohzfQnO2zcLEGTapm4Qsgozqu16BlzuVQ3v5Z86K07oy6BY0DTZywhymuGWvVAhdTtU
dvL94JKIotjkSRNJfZGk2UmQdF1Av/p0HEiW5wBwl33v++YKj3YAAxg02cnlGUOyFfeRSmz+1ctu
KHgJHsfGmt0OeWbE1iTV39nTLf5IijhwBzhL3xovp6Lf3Hwnf9Y1/9GZ7TWTfZj/QCiYPupSPwrK
rejMJOQQzFRdadO6CngXpM7wRI+LUek74QseGDDIHphNDRh5tlbnNQ1iQM6+3m9edMYkAZH9DfEF
WBmD+ilecCQjIbxPTDvurB3ohZ6kP88UOmwvTdOT9U4A9wgaKFVEJMC7njyMo/gGXg7+QzUt+xyI
y8WMf1Ne2s/OM73MBv5twNOjAQ9a30w38zTrS9u3qT06xNihYRy9AdxxdiPtFeRIn3sUZvrrAqiF
PwNcTzxALkOMLSx0h+vt5DGpw9adgCM77eSFkytqX+zEemL2AlLsJSwZdt5ThqNECvG5uNcvGV5Y
uo5OTOq6GOk8Mymga+DXlhXl9xu3g2pgbJihFjv60AITM+9Sk70LveILft1m/HLqO0i8JucYFcIf
eOzBKDS5usmYPK8BCmWYNWOxIZd0grMg8uCbrmB5yaQ7AFZbiLwdV4LTRVc/WFh/oUIcptzV2Z0I
NSEpKkyeRC2wWqdfEcGIWF+iBZDX8y2YvqbJIcb6RfKyrU9hEOd5wnbaFOUhO9sl+rQ86wlphh7T
IpnBcu6hluYD2jvZjnwud/bh1t+XiTHXYof55mEUUeApAYpCTfOxB37HWG07KtljKmPrmTma+aDu
VErn80HcW16AcRIiXpxKadYELsWExDzn5gmugfbQ4pItOJzzlJ12YWyPKVXqFezOn7u896tVeTnR
MX0RHp0vROdL4ERBjlyHmuUANat4A18CaXoBSa8Zt/JB/a1oseJ6ESxGSiuBhQ8NqSIO8WBP6lpN
Kdtxf1aeG5C2uyoyizy84aeISSxuA8VTqKMPvTq6mAqg1iRF4vN3hS/knmFywQjW9TZVWO6RO3Mi
o3w/pucvX3L7hb8CsSZpD75Sli0fySWniaf+nm1087Sq7Ho6IjRZ+lBbJi9QIZdsrkS1c/MNUTTG
m1nCwrG+7UUfA7TPP6vkQeCfU9RnJhD57rGifoJ5ENXVpvw0q8h4yHrYVVyUIMf0wy4MHevDer0i
fgKqAINVkIGVDtxCw95SAgxhb++663LW64a4vZHmrKrIqLhokrRcxvnuWePvcNd7hG1smxblXBO4
KK5n4ywWsMW8NIG/aP0T3heEtPKjt1PsaIFHlB8ZQJCYK4jFLSMZm+XnMqxFhkUUI5vIRf0JKW3n
7OSu6kawDPh3hjFgi4P2gxGe6FgVpbiDAUMSzog4klLgS73G4CThjiSxLbRAlw7I72OxMLjt8nA3
JM5FbffqGm1m/4z9uIe4ZsHk3Ow0pqKlUG6jK7VNqDHRqojAltA9PQ/XMI9VWSNa9nYj3iSbzPJX
rOLSAPHiC+8xrAhFBT+6//0kPYsQUaI4NY4jrcPOIK3hkGyFPSeoKoq5bmmxaCAI3BkY6roGIrJD
K9hYZInWuVGil7Rdf/vRHKi7pM4KVZ7NPpeb8WHMhFfcsrpT0cxpeDTV/F58/WisBnJqllYWnnX3
uSgNvx5wgz9VvFnYeciZfIFVBrLMK3B+gN6qq8v3WtmLHvs+14U8DUJHXImorxatu6g4wyb0EKq6
KMHKnks+HkKpmj/as6TIWevNpndXpIEPtVnZqLir3+KYWZC/+OCMtwnIsW3sXMy6XbjXKcP2qahO
p4VgyZDQm2zYiXacwdDXLlREeTFaau9LxTcENVCeDvJU0ispX5MkMe+Mrw5Z2p7YhYeF/UKEmBAm
D2i+eqJJRvVh7XP+UgZJfPGeANF7C19mkXeXFUlE30uuETqbL2hCZDa4dte/WGpujwzktaii9Vzf
Ec0qf3sYe1SHAIcgFcVziqM+RZ5WulvgZGS05l/fIn/V4B+Zhb1n0FoFIepXBRsnV5g1eV+lkU5I
XXR1MI/yaMeidAB7Zwiv+R/Zf1Zy36CPGdcEfMuy4eXlGcBt1UDpoR6Uw4lr2IGW0sOYNZgj65pG
5Igw/JS8i+6sLrgE8Iblo9DLNE8sQZy1wItzgGWQsa9MOv8kG4xVzHm1FJA22lR6xeKjjAPdzzA1
nx81BS0fiIVZLgTL5SSy7BF9eEei6L9/3o9DPHD+A2T8wqvMsx+wUDJsCES4g8Ug/hLA8O6aXAZS
W0PYdaIQvIiDGbVkWMudPxplKYkgLVdSAG1Lp6dRVnT4KMut8FtID59lfBLBZI+Cwvjc/dWxtU8y
QDh+9PZiMCm6nbQKwoZlXRrWA+yLf1pM9D/v+mbNBVJArxXdUM+L6GH9WVSPYkE8n79vk+SanNFE
WS8Pu9tMl/PdI/9BfBpe7TWtUVONZ3kngkQdaV+ZWui/4LyXsZpMsdsqmzgwSZ2d4O2VTZugv9Tv
LgYsbSmLBwHMtfqrDFhVjfpGEdiI7t8iwkwvAagyZkHtrUxh2yGO1eEPXHfoKClwnCdYEyjO3xU+
5sHzoDGYXK3XOikyu8U/mwsQpWL9ycheCcVycCjYmDsf96R/upftuQDaI9ZjwvIYRids+8Vmbh7b
FJrdmAeXhLotUBUA6Gh8QadP+obbuesyo6Jci+B4SlykniwAhsr8JtRsr1aDovSx6QXx/pIdQCC3
gvYcqYlXV7YdP4k8PkmkgkfJOoxt5TRg4KTu6BTiUoUcn42vXlEsDWz+e4FUx8t2XpndCFlTZJnP
AViQYEl8skr6QFE8itRJkB2ClGKP81tPIUNt/0POSvEvCLukHhZfMvUJPrzjps0nf3nvqqO9hYcM
Dbgxunol+ePi3urNegYJNV+0y0nhBxIwNTGY0gXJiONzRDfpEn9Dh9GAVoG9sgLbHM+NwOEOQrlO
yQ6ziIWu3frVqP1GBqau9UdAdugcnQ965f9eI/ijBBRRigXTIeP4Ilx61k4Vx6yBKIP9CxVM9K7J
bcFeM9CXe2G8x5qJ5RTL5YK9vvimmP5TjdyLCvhfv2jHHexQ53dEUKHcCVb3mV99prEO5zJfyQOJ
scTjBGBuaoeAZXDVi3VvWSILkbusPMjaCWSs/TzlxzLE9DQr6vPXZH7Gg3c7Rstsw6jht/5SvCQy
W7FwNXcCkhaty6csCuvQDWHYc5Whjp8zEUvypnC1nJPQh07o1JmY+uuYLd+5UCiUsNNVwsvP8McN
vVDwK0wRl9/CEk333Z2UgCPH76layZsJisnrPS7fIeUTVuj8xtjNZl9Z2MvcI9+HLwVvghLngErQ
A6D2Ma4/Xdw7HVGQsWiLAJ5V2fzcsv3HJJobR9ZKxGFx076nCphlyJzfqf5FQac7gA0WN+4rEqJr
YnV7SjC5b9mUUV8gbCEYbeqgmbc7l7AmoaTekd2IBAQg3YBtdc2Yw3KPhExMPiIjpgitVZ7ylC7F
A9V6rF3mzjuUwckavgIDS6mBxqzhTL5WERt+EOzgyqwy616NYTsukiXZ4ssN5AhbB6K2Pz5lC/Ag
pf+9nv62MoHRvCR0TovEjVwmC8rKfVikxHWivWel95u4pZrLzknhulikPEVta3aiJVje8SIvx2Ko
RWonj0gRg+GTG86LpI24TFcSbZkVB3Y0p5F0MTiGAgIIEDouEq2u6/JZiX86/wNXoJLtRhGbCD8l
tx9anP3PuufX9gJaCMF10W+XvTkvlT0Cw1Efqlpt5hcox2YgPuJE/QJB6UQQzGeJPEY9O2gXB3aW
TjYZpEL/HKejvLJGJZHRmvuYuO8d4ib3OodmsANU7nhplpm1q1KX/iOc82ec9YkpKrx21VY1gNQO
3KYbanA7RaUeTLPvR4HdRgUvIwFnsDKaoT0r04s2W57UAkD3DvdrQDDrr2mIF85Dafg8b/4dt9ee
8odDI1UijECWhpJ+AGZSD1dovQPENSDcW+dflWR5t2U2r/iwXaKwtpc9H2GpoQ8Oy5AKddNLPy8r
mgG6JJk57ReNhcA0IxsE8WwZj4PNOn+xol9o7IqlOqhtx7zsKfLXQDIsTSGjEw5FrX85c1Cul0CF
ILBwK8j/dbXtrWwzXUtHc2Xg2c2gdzKHf1hS0snvjt4IcEq+mRmKmyS6CQwLAZJWxmbMCn6qdN33
Y3jT93/3r8S0rw8F0L45zhfAe/pMXJli3a00dyUS7RYU9q3mFSMC04DxapHmvh67ECfea5cMlIL9
w2yCkF+719+WI3+kqYT+nKCD4QUabLXp67QuQXUCJ/F+FP58q809rp9kqL5bikVVwxkpIwjWOX5b
Toz9IhYaFJJ87el3bcGSKmIAZ4fsY3GdJUvDzyofAPRPOQRXLtVPB8u3NV2DTGReCgSZ5WA6xGJM
mzbQmhq3yXEl79TXHTUsaIQ8Je0QjBIrOjHSISaWMXdlace2G0bxkv3b2gmNnWwJiH4TJEJnkGdT
lBD2UViHX1on37J4IJ38niKZyeD1Z4ddKZJ+Awgg2L//wR3eQTbPTZNIFrqbRTdo+cM/4JSMyZR2
9Dc3UtM/yib/tpCNvBP6gJv9LzI8YvkkM0zu8jDXFlQ5hz92jAU6Om/dQ/RPyCmD2CXZhL2S6bm8
h5i2JsZGDiPVkIfzKImE/AK0P4JyW9M96B5PNKHQV1ga7zARy3KN2jWvXTYCIMq7WJ9Ehx68TApS
rzw1KMI/HgEnoi3rOJ/fCjAVudE3XvoDSvhD/U904/yhOe112ZQXY+/yaae4Jt9i1ldCZn9hH92v
5ED9bBQ5nlM6xBjyLsDMVL06y2muctpUXdayi+zP8jQ5kHc8/B8RqbfTueIiBhe9JP8vPurxL21+
8Amn7dge8Uy37VDPYLClEMabcoteHKK5YVxcCjggMfkw/pmJpx2wmN/+0PlteaqPcw3IlQ+ihHyX
2aOUI8BVeiPJtIYOWHTApZIxJmOGV9vpybTZuM1T6bntw+XvvJTFkpPRPP5//7JeT0PxJNYRsNQ8
4/GXpt1wy0k8Phq4GiJPo9jOXC1c7Td/+nd6bVtjqi+ScxBvk9gL6r/kNuun4GqNYQc+5I/rdzWx
P+4y1EhEkkJseHfE+2H7Nyq99pAt2IWVvVdcjo7uxxkcWl67kIVhydGSTZQHwsIYnGcnDPGh9ybf
1+VddcCkGUsHDodMFI+ftONuNuOEsez1j+munh12yTAAiRmE42Qt93iAh7h30+IJ9ZchXpFLwDBz
CSGW9jc9iigI3MI++EAqowCrivRuGuwoSf+IOIV56mYePqcHME/YFJTIQxzTx19w2JTU1x8rIaXK
HEKBomucPkxUXnaQySozMbe13kgHBh1SFNxU8eOT1O1lX/sC2yfpxpPGCQKNi/bwOBCo/GRqCfuP
uqwg1jUIMgbOCxRSWfqC2hiVZIWXuKOFiAK8BTYdCUHBAyzJXhjThGoOLjfjut1xOYQpZ5WLLPGA
QYzNX8wlo0E+21ak0WO11JgG8A3h3yrmZJ1TnBC7kP2osAHz50htpM+QeNga3tHP1l8krPrCqZ4q
5FYWoZjt57zY8zr1H+OYrOmlN8xmmIHyn1oD/C71ZU3tseGqudBw6RaKamvOb7O3twScykM5clle
XqyalHrXseuiMzS6YZOv0heC1r5pMrKRQen3VoyY1DcPE+ZLaF1lvM7v99z65mOTvgf2Mkp+YTMF
GWzIAJJg6aNgj0E7U2+iWo/odWCvp3J4m8Mk7QUO23HeV9tfil0xOZvjLjTOu8nU8RItXji6SE76
ecCkNXenYy+m7GzvHDRGLd/ruCR942hCgawuvKfB3l4Oi9jI+o5iRAKojJdSMypNlNSZNEsk68bx
YiQbFw0grSEUJloBKsgWCzTwD92P7yHi8hqf8qnRalxM4mHMbLUvuetA4TFEs6oppGX+qLCzWSZr
QRCZkTtemgjpp5Dlt1ID1rdSh98rNsDz4QluhDy8piyNemtfGmGPXFVjmxF7RmqPDjNIp4dR7Jje
tBTKEsShbyXzhECs2IlL7P/3WMr0ctkYMpU1gtySF0vtVBTGW3aA7oPYUg59J/WQ12s7YNx0GwRl
86hV7eQSxIYmY9wezOVBKngfDLsHMC04YJoDEwzg3J7HGFXAlQNrw/eMNEeK02Z3ZyZp54dEubYs
cq2zJqnZrBzfPX6ws7XLAmV01O8T1yIGfP6MIXEVsOr9+Gn8xlt4Ace3OvYnDQzl4vnbC86KvcRf
GCsKsbyAeUkIPqEUkPfM5DFVSYdYO412ot5gn8hXUgeGhGXgxW1To735pnhgz/MF8mbfbbP/UCz/
AMllmkIgLM3NKkDHpZWJO2x+rfJEU0rnaBt2VwzyE9PsDOQ6/cgakE+uqMtTL8ltNxlnGfa/CxQe
MU6AZM3RNPDoBTIXZsybm8Ec2tuEcHSNXrFD0r+bVj/W+uMA8/HaqcyhUoXLUq+PLwh5sUJvApso
Md3tHrmvBHCH1IrAU+LmR5LEul8KZNysLJLBZnmiWLKsvl7nm9ZnTVd9O3r4fgokYz+3VSMZgtVB
Aji3MclNIHGnvHuh1iLUhqeVc68DgMkkGYySIjSNZqFAneXxVICJ6/RlH83BiKZte4A4nwe5P7rh
SDhf7v+v1XVQe1oOb5cQsenUn/N4ZulyxoXGa509rr4Qk3HuIyA3M53Nq9D2bggEhAbJ5/LhAFZ4
do4CM8a21DP/Ko7pxQCbWyCf9+v9X0Aint1Heo7wUSXNJS1+2c5L20M8B3JrFEJyFeI9YUxCQ9Mr
98kNffFV9vaROLefndRsRzwqveJm09XUiRf0EPn4PtPY9bkcppKsYFhJS6HQqsP0qBqg8ohOS6op
dDkbdUnR134P/yTbpm1PJqjZmy2x+/GHUAe+E9EWn5vGdcjB9s7MdWH5miWcQuLqHmH0UXHsqHQR
RxgsVyaEINNXWdGSgFOXeKXS3UgBbu02WP1Rg0947yiq9NRNjKAcgoxMqy+xZEkntnlQ2jmNuJ02
4um8zkqPmIXSZbdsRvclMWwuuP8TMtWP4WVfARh7I4HQC5XPCbTZjKJBLM08/ySPE5SEsTMHtEub
kssloeCZMjiWloYHMvGjB0S1+oN32/QqJbnqsgYwJEcp0cRsBBJhqavlITc/LFOTv5uNPL4EtBhl
blwZVlNf/F4TYQaqEPDn8IXYZmhOI7EmOIFpzGbtdOUyO2hSTmA+gUIePZQuUwpkhh9tijTKkHm8
e+uPZy/JAyIxdyhlU5ynUd3kNRAfIrOz+plJTbw/+R/GOcycQnHsbJ61aAYR3dIvzyeZMEeUZQbj
RN0lCaSJb1ucRMiLwlaFTC4xdPllKVOYmUaq7nhx9nYLk1zEYqXhcb0ZzZPmnclAEP1Ize3omzNw
f3P+/zwUUQIEPeup1WxY9x/CPjy9mgDrhMmIPRmc8tmu7vV57cgTRJVGwqh/wAGzassmc/DTMtRA
TBH2oHpKr6N3QT88O5BBy9Y4tTV15NpH0cZgLwHgdwtNT2+7OMJtrwKgSteiAMsVIJRFsjzqDJvc
1t3lsdqmSsRHnFeqDBgipsOvsRtGiHA/wWb8vrAMu9d2JeEO75oRjht4nJXogZDZLMGwu8Ydet6z
qMHFhgriKiRykItIIhZmsjggB2wAo0lWsrf/xytdFfLcwNK0QnT1atjmM7/x6KgcPETEme+jOvdZ
wH+9Dvbrl59a2cjd9k+TWKYsI+C/G3ysshes13AUK6tAR3jBebYnejXHoEcFC+JLQzW9RC0Kogul
iX1njNQYeaoW7nrPEZS7/2ldEqYGhDCPCalAqxDRINzorg/dCTnQa5vc2+pADSnWkFIb69ZQK9r0
D3J4iE7tmqhr1JmD3VM5NimcBd1hO2CKSZI/KRLLiCLRMDvalhdgnoEuYVZDCRYPEYTET6SrROce
cmNqRf+NpGjVCcXRKxXGeVV7jPnedvBGF5DzYKkeQPyoFpRX6JgS3o6HbfqqDJqWj3YbDRb4Xm3+
yy/0FODicgDJY5AqoAW6nr3mkTRyCq+ohyTCs35QWpR+5Kv9jAlPH5wEDtXZbxXc7QSJWS/wnFCy
Yn7X42MIlBnAZTVp+YVRElfph87GFkvzDRnFFTEyiPlYPhTWohCrFS+P2OMp8BfbzvgBgLbOr9SQ
9p6H6MgKN4DDgz8MMfWrMspGBMieUmat0EikQnnjIff5uSZpqSkGgf+RSkH5c14Mks1YmjDoo74c
uniJH0etwgMoMassJox76on1o8f/bmro+w3E620VRXMcRnC49/aRn8U3VSI6oRO+6aetZH68DZJ0
1+hRX0rZFa/LLhrAxCJm9u7FVGEp4B0IOLUKgFzIZm59F3uImXz+S0a4K8gsjQTJByzUg11f/7JN
6VnT2ZAZcpLNzmCzAwTL26V5KXsjrATB4YZsq+kVyJLdfOtyspaREpY2/lb3gb7irSCaMFWCjv6Q
Hd+HqyfTAR9cuOEvT3PiYhFZUkdhxKmcWSV1Cx9bbHq0t2JybOBdcgdmXACma6kPQIhfNCiVXzaU
a7O3ESR8jqzuew47LomabmcQIFh/zbACq5ODH6KAoye+s4qhN7UJj36441F/cVEYxyTdMFBhfv8s
/ujIoGvHRZHAFLR+Ug77HoMI8Hh4bJIaLABzliEmB05GKlSv4zBRnwP4rHOxZpAx/iGmme4mq34i
9yAAKVPZjYNjxEMBb2QjFWCCAh42eCi9vCZtiuF+rN3o+rwhLI+PoPludqbUSog/nI6B+KHHobOZ
gfOJnpA7bM2pqZ+Rls45D6APXoWO7dABuyRaxjL5y7AVXQ0Pw6GKrMq+Bn58mTPopBBglFp3ScrK
esUmn/EJlCrVcFChFIKd0UoKRXrSttm0ltjbpcXtYRdxwy6tHK749lL3yHw7tulecrcFsErU3DzR
3X/TbaUDPqPMaVShVb3OEQrknrwycxXe/BxobtIaTvz/6Js+fxUGK9ahwQgR7k4nyALn/s0TmuCb
fgr+JIEqWBAIVpn53jcPnb5fv+0NmMSTQRdCieH9MPUOq0d0Ulup91pUzL+Acfar6WU4VCaw25fG
lUEwepFTBz2eO5m/iMQ9YRz2r35R4uu9bOKaN+SC9tHoqjiShieN5JgI+sIn+Hf4YVNXXd4htr+U
zBCJNjdtrOMV9n0GlU/RKVRifM0lYVRbRYMmMHC2yQYH/eSWSJG40zF9HpdXN1ssoVxc0jKF5iUj
qQydtflhAXt9QaeUZmlX9fPi41WWmdZOL7pFs3ZZHRe8WzDDqOrrKqnAWrWVkcQuZhKBfb1tyz6j
+2DZULc6gIdO2rvRYmeylkvS+qn82jl+i5JT45i2Xh13/Ho2yFti3dlcly5hR1V3HX29cfRE5bjs
V9wbhW9TpR/7q3rAvACvBoedaWMKKHnJtRd4jPFgM72IwcNyCLL3eQcT8/TfAHDXbpj2BQ2RgLTj
pioPU9gCGKmmXHo2Dgmf43AXOFHN/G5P/rrCLk+OEplyCg6S5vrxGKYIxQo8m2hivlHE37yDOOxb
24+/+3ndXOO6lEUdG5f9m9V11Zx+aGQ6rLS+f0rWgGzm7e//Ih9nr9+k/7oEnpnYw/itRcmm7yiK
9dcoQgQoxGj10kT0Mdaf36ehJLb1Z4iadOeuxSd7peJzPaiDKj4Taw9iQRo1WaMilpYcG7dD+Hgs
kz3YiDsUAbgVYuOATFZdD/tR3Xnsr1L/4nHjVJFHg3DnMAsjSzgO/vbCa7vnCPhdk9XSVwNf0GnO
+ra1gm85ZOtJPcEjVrqDNm5R3Vp6kJ5GJe6IBmPRn6TyAPkobDRlfkYxw/+BQZkAbXTy+AZEDC2k
QPgH6QCJB9TbcA9IwO3NHpLGAX8UpfibmlshqCuDboQ61j30lKqxb1MKM6FsUuuS1FbiFI51P/Kr
+GlWdAT1MgQ+Bx8FT2mm8eHZbO9aXAjSq/Gacb03pFrWotdnm6HsN3k7Gy7F3avCNaG8QS0O1K4d
pvV/Jtg5JJmpGeoF2datMeBV+618jqJvqG31VGzU3u89YqjQPUElFXVAkM1nDr9x4sKHfh1U8gUp
jKzb3+yu0jsLtmbOW4CAPnZrxBJJvYCOCD2PptFT4IstRxKv7ZCdEiG2lJI5tf5wVoMkvpVPTb0r
u0tnDimQ5DTetLfEokGMJAxuf4AaTTXqErSrqaeBQ5PEOsOPc54IovFZebdR8c6gfsRiwrvlVZnu
KC12OVONET1oRh/k1nZPaiT94Nx7jtozx/DT9AQ8tR77qoM3Oq3zPdA6h9BN5JQRxhePAG5G1laJ
Qdz420ncLRF8L/FrrjmZ2yzZFqI55txPnbIOpbPH5f86ASikGGmVrLbW4eZBSsVXlDs40LvpRErX
Mmtf7haYVHcB/JRFt1p5fHS7V2q10JaZcoXRWlj/hjSKQ7ryN2EOHBV2vdLLLQ2Us4dy+v7lgFB1
tmEO/SjfkAje5hLC3nVbPlJDaXmrXOPyCx9pOpMPkfRR6f+P5QOX6PKBf10SXZqbpUnKTxNb/ylZ
sgIIs8IHUZTU6ouWRCtIx9n7+DFta5l0mfgZ2FKvXU+XluonzG+OElTUwG2ObMdB4n1kPePUCPQl
XCTUoY2fQKNHCyICjhcT+0PKWVe8C7kPG5Twd307r/zc2xI4TFfI5oKCPHg+rqDMrHBJYOzKCgYQ
KbS3ZMiTv8tvo6GwyYE28SP7D9jWVSERoqpIFS8UqI8Ir8tZqy2/iFYvxbHeLsdQLQsdSpn7roKr
6Hl+82JdsYBCjREGbITCQDIxzNRSQc/VRTIs1jXWtLZzeH8hcGoMPah2LjNwRwLQY1A/OSkfIEPS
lZOlfj/qIJfIKaTSpdwVhem6rnnA8wioeBku3bEV5Vc4WeImk1nuv+lk7mX0t6ASvK9Opifwx7AE
gi/WwUm3e8KIlIroOkAEg1/S0zcq5HRaUISk8sJMpmRinUx3/uVbk+lhKsvwcEveic6ZfWLhUhjL
Cgu5lRpCrwhw9hF1ttMdNTbyiEdq3Lr7YqQ/FK8dVJ/DsTg742Z4J56+1V7UkMsbAiPCdkfZxv4J
/6syKw2Yg5bQdHhvda9EjUqB50ubIWOs3EXbpMZOgwOFmBth7KZEqfx6f5x6APiEkKBqiSpQRt16
i/P8OYdLl3cUiQdjhAv56eqZQgt2M4Ide1dlFUjc2ZVyY4pXpSIZ5z+d1yt4P5uMKYkwrZDcZ7I7
FYTR+4b5J3vFcsl6Qk+HU2VXKTWnbVqu4oyaPq/HSgVuVGW09cmE5yJtH3SvtCi/kePbxI7kcOQ0
hVVGFd/6Rj9rxbc1ohXBbHSMUg5ZxZjGyRhjk9Wprih3LDpjHJAZ15O+HBEP4HFio77VBbObus+R
t67IUZRrsJpnWajz+v+vFy/Fa+774J7r4yQK7K6iM6QyB9yPRsYtwDY4TqU42jiev2KFVUb6l9/m
+lXVK9pmmtSUASeIIC3totYd0VumqmwXCwScWMUVdlDKYOSc9uh7Rrkeu9EqFRMphBtxI/2Iwj1N
0e/4V/knf+oo6sjPStC0LvnLJhTEpo/RauVNQ2xxqpnCbe3t4qh14ZKgHxENT1ozjqHYgvyleFJW
d8vGia4Jzy1JZY5ccG04Bqy/NAkMH/m601MzNqfjtvUgiIE4O6IRfe1P21zozE1fn2VuG7MZQLYr
AGUpfJe3NdXVW399tgbYkqiBc9lQW0vjndzy2Q/U09MRd0a5CpdJTzISzITttXNDvXBoTbShSAYq
cT8wVcKU7KoiEtrgf8FrTISYc8XeTbWhRoPlCT82OoRC1TlI3eJ44QdFm1DkYAZ3WNG/2dFa7Gf+
igYcp0w9xSG/EqMyJzT5bS9Ah5DtnW77rFJA/kgHKJU7XG//3w5mHQNpUiGfqvQbr/codl4Jzm2Y
1Zce/nX1plRJMRgZQ4EZ1x7BdCUEMCYPaoEvQ6C9SJygFuev75GWKVh+5j1891bGmriZ+/nDTOsL
K4eztGP+egoNAzE9GtWw8lMPE3yBr8U4qUF2129MN2vTlTYXNdx2ACyfZr7RAFIstmuutEFziBm8
vEpbzPUVpyDXEmJp4clANUgVVC1pcXlczSa7zf4RQBneWSY+ZpdEhf/vDq4lu/PgLUsiRi7z/lZu
oGFdhqC/3mIkD9WJR24WP6eK6t5gQacEVTrUVs+9ZHTH2rqqIxdoCOCVKaNmcSBMopmKZ23RDS5v
pSZGAyJfwIKHLlpnAhKICS35ZuJ2xDxgHCfao8AYWvl3demxuc/HimRcLFN19UKok4kNtpBz+1M5
Z/pozRcZPupadd9t7ejAgFSqCszuRNHQC796Co+Ix4/+c1wc3qQpGEe/aj0F6v+fXgTQg9IHRh26
Ch3AaBGyx85If3v5P/7sS39cn+MgwAIom4EFanY9lfYD9EsX/vEvrqWAs7HQP0Sp4gTYjEmwPeRg
WyLUtGlYkJmiE6nbxRq3JT5UTR2kkmnjXwS2ELtD90c12vPKLfpi8mfdIdHCiUFdNlL460b7bRjR
opaqZ62JsmuwjEuEf6cpsrSV4Z6irzAtuEXE06EPtluAtXwknGfe+4vrBmQbSpvGoSlPUdnd1N3k
R4XL4QAlMSvxDcUjEy3HOzfSBZXVYsWbEKnRxe4ZRo2Y6186Yf4xb4hBMhgF4rVii5LgiDR1FdBY
AG0sSQe1HyGEDewxnNwCM1a1A+bDVN1kvzJdm08ykZEQwbNJELsXeeWplNDf7uJq5931fHWxqFCb
wS0x0fWPtD7MwzMtsXEQ4K1xVrHt02naI42nLdNpjOpK+VXx2GOztsnogQ8LJ7Wm8kd1GNR0Bqls
sV5w7NbJshYhgRBU1z38dggVlAvu8VU0orweZK6ezzUYNYWBWlgIJiqGlJ9HMx1W4INPFOLYcXpP
mdKX1LMgFmQpu9CC4jIbE7zgpV+4sw36NtpcugLA0hCtbBQPJtFUxSqaaDyd4TFpoWwf2UnFyqBp
E0+zzgljONaIG4BeNjyI0+N1KKWTYwN3zFdiICYlQdrzyQNa3AzkwGoEGDksPw8UH6WjRe7fDB5K
DnXEfUfKUzBAdaSSX332X9KStz81O4Fy2PG8MI3MXDx2yV5Y0ohNUv325HAw+t7IqO8LR+Eha533
jRroJrHybfmB0G7u/zuNVTIORUs01bh+AjlV8mPhExERUP/c9GxveWRtKpnai2HaIE7DQrbxXV7q
OazYH6f9QqlSTT/HvnQVs6CuCNx2zJ0oCFIaB8dE3NIkmYpxsD+p5XgBURSIgbHipoqEpIAtBnDU
X/NByiHIvWkkRtfur5SAT5mrhM5j+zLbsbts5RSbuFKSVTKwt2tPk08lUo2nxRQYjjCUj0K+Tqqw
UQe0JY+e7Ctlb4gv1N6OlPYCk1ZQqo6IvhxS/22XqyP4czQciF7c6Jku6nFlSBXhm1tn9k/loXEa
2ruwSR69XzI4fW+Dj2oNfu99xVSVLL88Bj3B0TzqtB8CnJbfaOTj9ln9V1SJxUEZl1o/NTkLjDoF
fXrNs1wPT/Wu08dAywGcm13sfpG+zcWaWFwaP6VfPmHoyzImOK1DQie0xUZzpEyEoiMv2i5Ul3eq
qQLUpG1xfnu8nK4egZYw2/Pc040bDXjsullgu7zGQXFMCcs9tSSJEyKlzPeSix5dDe/Gq0/oybJg
1uS35OYz2zpVuMkL2tfDHNKoatCkXTwxdQplAL+eFVJwCQlrge20SGHIwGrbzB84r7w1urq1/QXN
pzgppYWQbEP4Y7RTuG59WZKjnL8jCzhZoJqF+Dugt3mnrp0lOIuMzM39U4sGvJuZoKg9evef7iCM
M6TnwBYW3u9OA9fxswsnnxZ7XbMoEOfynQXZUAYz41SgErQoDzyy52jo4yZyLnr+5cK14Ga8i6Us
5etCW0eJTvUTiOUuz63Wce/pOqWRW55oucOQR7iodFmTfDNBVpY3BahSRbVKAK++nvUvPdziZJMY
EvipuvoAfTRlYyc4mDBkmaeMVoZAL4mRJES6JaXVda4Ro4cAWl6pAHRVO4u21YFJJvlUr1iW56Q5
sXQUoS9eU+uYwDChGMmYKxrkw9Hp0CVxbrOVhjSw4aeJlal8QAcE4+0ezFK6U/YM/ykU4DydFZgS
4NUTpKZovPM7i6kwrVbhR2mOuGk+FXcRrGAThV3/eMA8/coj9X3rbSx8ky6U2HEBNUUQZ883vWxE
Ee5NP5VK68t/mQQY3S7Itn/hZmnmRQo6Ns6h/EWgIKxZS43y3vHrqpmz1CVCGgtT9j5tH3wiRf89
jAs0s/6yPZ/F+RNhl7jtRRjNP3itx8tQsxtYLAXjppwX978dy3aF4bL0YZ67yIFBToJ5DZk/7mwo
PnNFDyioM8opUJuzrktxeRSzeTaSzWSDdRVho3YyO9/sINCk6pKEZWzkvkezA0MSDEiBtCCSGWvy
Oy4lp6XgC0HCSTkCNsmDIootetPT2gqfFATpWJzsyPI5ilF6kA5uCV16QOTbkXuVhSZgVp4sUK5n
Xw+8gOa0itA1ljLxCULfJx37cBN2zs5T8gGGk51CjkPQhuIvbRn4PyYi+muEGMOtuEwP5rcbnmWb
WqEfOZWrvgzImtMWGSj8fze33ZKW3lvFcjvLJ1TlYhImWuA8NVByQCosQWd3PeeNz/bAgGps+1MQ
IkYcabjqNCce83TSSDNOvoxCbCVSUeJRYPirr3FkudOECIICvugKdEcrUzDw+wbpWQs8y51ei/T9
QHkjKoLR5WVLPvB8N4W15p0YzkW7Dz6XaS3MjOltk9Bu0Rqq19mmvNwxwXF3WrgOW34gxMYWm2E2
2qGQCmEAQZMauEGMQzt0SvIvtKgNXzE+53i1W2thk0JGJ1dC+VkD69/JneSgu+Kr9I7kIo1bhizK
kO2uVXPmSZgpiVr+zB5k8oMV+RNYIuJPSpUAblbfVHX1w2dilRLH8kSU87MM4Qjprpgxz+A8D6JF
fmwVjJJvGNk+mDzZx7JUmdgnM6BKff9tGLu3zrlGUc4GyNmWMrz1TFuUQjwcgSD6Mw6gusaHmLfY
a9oBGLQD5JHPXqdX8KFl7R63LyPtnywPvVaUKIKAeg2LrB4j9kFy750lVn/jenPLvrUymQSCwTV3
fYnvGtHsJ6uaIy0ET5siRRl1J0kYRK2Qomqlzu7dwr3cJjdlI1XVxJMHW5rRnGUJnMYAdp5iMSOU
gMXPDB8PHuDHTAtOOgWYq8pap+70InPKQcTu+iTek0N82WANkEw9BzWCbUCV+xAgL3rpejTP5RVO
NT5rxlHI13d/NgFeTFf1obhjGd087tLLD72YPDGSrZjexvAI+xTIHv4MHy+ecg3K+lPSNYpnVeOz
p4D6DnKNmYg61nJutWSKd6+8W+WmGoW5+C8w3xqeMq9Ex/uP06TxMn/MY1Km5xEpaCd/nHl8CCCb
k+vSC8MhyK9tOuvEnR6f81R1pSYh6Zvlt8n19lsRGedjF+O+h/Si0NcUTPsPNUirvJKwouU8p2LP
5PAFO6Na4vRkWYw+yz4N4dJ9MC3GOiaZ0+35DWrivrkgKci8UMgoiNEf1+g80sb+8J0aorkT9NXm
SO46y/q1PeIBmeZklCXMPNz8SY1bC6n6Qffqp8wGHg7xv13jfRUK8aaolXbWrPCOcxqMrvcguPwl
vAWq/DeH3lrwIr9+QNhIxOwRF9NxjXp2xGpnrh6YdUez6wcrnqrTOPPkVKSy87SBZCKdtwY8suhv
GVNqCofhQcrfnOb9RYjLJg5CpsIpfxNlAG8XWPIG0/H6KlPOeSgtPHCDIOCSIdiMXXwz4KTG+m1W
hQic/WrpAWMy56Xdc22VgtdOSTtygJL2O8HPx1RTQ41SsX0z+5gdsiPT64dNbI6yAnqN8zzjjsKK
B2oRL0K3B+BhdR265lneeikJj+pyBUJ0sEpHo8xcyIi4ZZd1lCjAtJMTmKG46lvtxiyK6PJoJ/Nz
N91YkJRZSXvWvOxZAorxF+qwhdsfJP9Qre+4CkzlKqRzgnmPCo/wXNhHAa8eyTpmob4cn1jeN8B6
WtPr+qTxt1wc6EcypwmIPy0hbXtZEo0O1sdQNUzrE7c0f8jfpqjoFe1OhDv4i+KCywG1zNRGNnJk
5usacimOEcDPrp2jPtflZYPjDkPZ8TWIw6Wbsnsm4VzCZMyHi+2V/++X0qQi/WBpguPqDMUoqCeJ
gKFIPmk2iz0XxcY51YP02CrQDuCCtHD7qN1Gzz1gEfvlu6ilJQz5CDNyU4C8hav3ekh9x7kI/47z
CWlGBg4N/uUo8UoqNfQDQCG1EGAqL9EkakQVGqy8mRCc5EyGwxFcd32ssyKc6GIkol+JoUkWFPG4
bClLVrdRMvfOoKT/zXNWVp3psDuzoQCpKvCoYoBD54lob6Eq9JDfzB+ZKGyjSbyJzRIEN5UsoCEn
xncoKpqjiAnVBAL6sLf1gJDWh3O88/KBQocbn6a3O8PAFfULcNAmzGDGWd8WYLYMxEu/hoZg41a+
WqFTNuJuJmaHBknDKvCuNROAGIe8gbqIS1KHMkI6ra20weooJPvU+ZGh/kcUzDwdVABtPfCRpVwb
3gTV8HaQCc/qIGGQoBlEnGh4M47rcPdBHaMUDGbwERxYJfYND8ReccKH0jKEjrNBdNrpPw9t+FaI
N8GCAGAvAZBKHSD+qcU7nBM/QCUuoY0suOTONpGFJb2JzZACJ6gtkAIDOrbrfPHpmsWCiAKxh0ND
zgXKDbkgeI+4qSDIimNAiqf+K+49cZ8tPFp8EAbAUIOZFksldw09hQ7rs9v89GFvMiS45AnlXwMF
6Kt5zP2uOW0049zv3v3UU++hoF90LjBeW8SCP2Noo9JBModWPH5fHJC6r9R2zjAZFw94im6NMHPq
xNR2p1XtUM3/d9XdZMXHwgIT1xdLaw/C+hID1waI/p+isHL+Wv9Crwyk5vLsSFQnR9h9T47DvuAg
ySJj1IMD1Ut9z74ITSU4MfpPh6+cHEj/9vRiy2auIuiL/t38/nA4m4CBm5CO0haJo45kHN6y6gwm
89uifANpQWeOnbMKcx0yt+F93JjW26Ref2giUqAmz5X9zomlHsvQr1il/CAiFr5XIGi5v7SodTzl
LGX/rldqg4RQygk4Rj+r1jD4phAMxQACvfRmdjzVYD6RRy8wLsAHqGC+wwjVHbTdft/dSiTzaUPV
kfy3AQ+xnRC1XyaHLDtjuGfDFoiE3+hBwkcmB0bEzVmW8N66/mE1Y69GDZ9NynWS7VhgfkzfU+Jk
pqjsRQGXW43qleX9kfMjTKyKdgh7l9sj1R46gxkPs/Gj+1vyuJ6VkX1yZC2D97tdHMOQso8uwGSb
ZySIpKXKLps7IxwSwp7+GNxN1PeaJkmAVKflCuOHEImzM6K4oiQ4uw/3AN+7fFmLXl9EG7IDNQx4
GC4strDBBIf97pOGKe6BIPYVHuzdHGqSRh5QuWfQngy7O1LMe5+qR3y9biK6zbtqNwZtx8WRdaiL
DiNlSuoJ63wu36kiMH6+BtICCmrNEymoxIPQjtPCkFhf/D5U1f+En2EQkb8f4PYFipRrSzSzirlJ
Nvhmf79H86nkoY9Udv6PuwHFcYaanE+w7vCYYedgCN77GlDD9NN/SzFt2ggXQu0K8IDHIQ76CnSF
BICGBI9PcXbInf0Zkz0MLbQumWdx6IV0LccWAL9GVGDntUHwvg4iAiwhBsJWYBiiSf/IK583iS6D
haMn3Usz/eOrUrX9liPV5e5xeQf5mNzzjg6ReHlYDV3GHEBSi7bjEY2KwWuHwmXlJaSct44Izs2q
deC6S3tvckFF1C0FswXUpPJ1ir77znTlQpxMNgYJPr7eLLWMtQE5Kg5rW/Mu0PwS9y6uzPIX/YYl
H5Xje0c/pX9hpgtL6O/+4Sh+xgkywWT0dq1c1JjviZxDN3iEBx6iaWeM9gld/1GLtIai0voTspOC
mrRiEVdseugmYza/Zo1KgFuNlr8bT88a/Sb0pKZ9gOEV/9FGKauvtoL6OxPELbb6ejLC1QwBrNCS
HL3d7YFHOF+2amJOalbkTNDY5ssXKMdzrUHGFvExws0e1hpBDfwkOWGCgWVHQe/qqUEJbNkqV3HL
KmppR1iLpxQFLPQSldr2fFpk04lY5oE5GeP9rduSdZ7oPWDCU3f06PW7XkuKz4rH603cT5NamuwL
IxltOBWXPw1343kc9SWrLpsKdm9LWvSyuV08LpbEnzYMBZJExXXkbWnzKonbDnAYbriMTEn0p8z7
JIxsR5wboBNVOWzkZ2OSTkKNimzqysKzli5BorIbPyr49pkGcTuUVRgXBfvBg5vi7WtqThAfjMdF
9FNk66NaNzqmerM+u5pMwsfEfiosdxxDWbUBZm/JEpfLMlMCi2ikHJ8WhIzCuiFRlFyoweRuOgkD
PpNtHjbVGkki+6qINseI5PaxtyVR48debgiNzaix8Ywh7iiFwca4E/BVjWwMvor6Azkn+vil7cqo
+WAi2ocKclDvSvpgo9GQK8tMYrfplnGY0MFvl1V/+O02eVoAyjZOw/2v0PFZciDVnLzGef/qcNQv
RLenwb4Yo2VedrhJn/COo8FazK72MfJ6OMzAsqTsTQXYuDnb849XfGD0ReZLIU5JhiiRnQMctxPE
uAD0rOlFRIgNAxH6xsrXuGuXROHan8JDthLrcFY600fLXN2M1YIDA4yg6X4JZzYN6N61c6e18YDi
lUR8Jg2FnlklKdtu0u2LXd98w5ykdDWc0yEzAjVlkKz27tkuWIWZdxtdppANKxl/AZFaxcqgjAaq
5qJ4r1SUiCzuyU9VDy9PhGnJX7AEF1oH984RUNTIbnjMFkBds+PXFQvo1LPJcPkx3OMUxdBK9+Rj
nwvIpLian0FGQavDkJ+Uj5uaOdztbwtVvdYvvJNQguWg4Ziv/C40Ajlp8dJA6Gzm6VkY8PLKL3xv
FQ1Hn2q9CES86jmkhYcE41TyyZ5kK2wSFwszY22k22arF92kvvOiw6LDg3Hdwvja1UNrfbDYxi0F
Ei4PJnPCP1oLAAizecD/cGNEujhMobx3DY5T+zK2RHPLLxBK/DCHccn2D0n2sR5d/lxRlqjEQ72X
QqllY/8i6ziC5FS3hPvp1crc6CqBlr3WLexrwb29KtbofhCx19th/YTCmSQ6tJOrS+VsXKtxCqIa
qU0r9PXjO48IH9d3Qi6MXzJtPLeL5j3P84qIhdRHhk1AkJDd210Vz/gEXY2vL58hEbSPATBcXsmQ
GcvNjcYHQP+rI7zjAW45I+0AWkSbxOtQYVA9YLH5spQY5pZSotS/NENpEnhcVfFnp3QrJzWFgcYn
YNkFfQajRIMdJiQzgjFwwXS7Phlsk4ZJqXnRw24T0vw4vsNMmc6tjL4WAmiYtUiV4kAMqrBY7hOS
vWczj6x7YLRn0hwZHqp5Ub53yPm5FoYrlPTuZK1LqNOq6RrgMV8+k+Todthvk3QfPfhtgbIzUvHB
K8zPlOLQ8RqLI7a/sP+mijbyk3b+/VpanDz1ru1YbfdQrgFH6Z7YI/nhPn+LmAuZcclkMxmYkERE
G+0FG+VOasgII0MPu9k0pkjdZmAHApnqQqdrA+YMJWOY1M/+OHkrBCxH/x+kbCy73LV8WyXz4pts
+3muGtCW/dmzg5O3Ok8amaSRCdgGnlKPhM+y85NFhbtEVQLcCmMqIgMIoncJj6a26aDkwv1eCHs9
IGDKv4hhKeDKltOaW6pQ/ODH6U8DMDoLxjFH9YqL2Uji2Q0Pg8Sb+lR1j2nkOE9gZaXakokO0btb
5mmLcIC407PR3HXBXIsWoOS30MLXqUOoUJbp5iPA7uJ2D3v6myHG1oV3pov3Tz54gpRa1MxvReeg
XekF69zu1JlSLDVvLuWHfyGM9A8gT0DwrrmPzDnNwpOJ9T6adSiHFxjqUjqudFUj2ibOsFkJKfr7
RLHjCelks4NfqmVmGT+iV5DgBVr22NjGPHgc9buvIMLEopbnRgIoCWtRxJKiQw3898sVRnFxVSm7
CcAyDIDyKTKhuYQKzBs2CBexprmKe5lDihJJY75bGSP29oakhI/jcPSP9Tv3C9W/JuRy+cE3PkWg
naezUePUiAssHPKv2qMxizjx9Uy/HFCfqkhGFcRl3RGKluTuSh1uevosI6ZaxF7J4uHyCvhHwwkG
JSysLd7Kue0BTu7+PERx9jj8edTMWavWKz8ZBpwcm0RPxZo1456IwXyxhaGyL9yj+S6CGrOPkHmy
ci8sfp7x/Alzm7+CCU74KNYldsOMvzj1dVJppochp87egL1TGgZ2SRzlDM7GnDVDt9GR28/3FFve
6fTwDKQ92J/pEFoN8zoiYra61J8P7gOZYrXxe/BYox8F7UCDdVXMzTI/Xy1IIOFeyIW/6lM+DFcc
9mCQBti9bbj2U6BQGExni2VnZUaKUvKX8pfcp0MHv+poZLHGu6zEyOObcav6y4U9Kgb6HpKDCghg
c1pkZlqHR5BKOrj81b2rYd8zFAYZmI1odaRJGOhvV369MSavB0OY7bQ4SdVj4TfwNHQPb/RYIt91
vW/KL91zGseJJaLa7faM8bhzJVGPRdL4MRMEOmBASwB1RwPZZeST+PTUHUI/xFeDHqFHBHMn79Ex
kiKB2yPkgsDm2XJ+bCxqca8l8yu8HGQeeoJklpSgqGHqiMVRQuKdInl3rPOhCDbWiUX9iPQ2jfws
0hKvizt9ZMmMduUMsjKV3A0mPGi90AN9gBKqEPnit6B6zCso1GIrp0/f0H/juD0kUcF7/d3yzcTG
kxDOKYdIJHJKfJpmqro88//r/8/2AkdqqGeE9gPxSwUmrwd06JHGgAvQD4BI01l1JbJcA28tvj96
ySZxMZ+D4jxtnPzc7S8kVvrtC00Ov2YspZc9U4RgmkEGbIQbzNAYSG1QVazI2zcTyEXVTmZRNvpr
7wsc9ml14ydZaKMYxX+BBImKphWnMUsP+HzOFW13KWz16uifpji+Z5e0XU1wHmILB5C2XAA+spa+
ey+zgJe7FWZdqTDAdj3N4t9XNTyari8ESM4Q7I+T+xTDTYJGHBfGn0GDOSVt+FaHy6p6tJsdCghV
jUJNrsOVT6c2QynOhnP268HsD9ZnuiWqZ9o8zBA7MMEtCVIQ/rEVYHG8ndP16tcg6P2D+srHXMQY
QwzA6sCrMNC0P85V0rLiEcuwrQ5+v1Fg2OxQzhU09XlisB+grUOKjDrTmyKuszu1pvW6FZFjK6/a
lBNhAdThddtV7/NJ/h928UQNrd6srMC069BUBratMeCfHNV8/qAMuVPHwJ5S+rIWC62iG6JRYeYH
Rltit9gVKeUt92uGuHnlGqiEivTFcRZIkAbqr3gV+YSb3w3aTOoM3l1dwysP03x1qhAf2wf83FO9
nCLfR3zNPwnyJ0Im8ZXQEkdaIfnhmcQyegGtF2uPX5eco7vZs59EGbIsQiAmP1IU8twQOuI/7AaC
tOJ6roZxsat95QFiWi5JT4s8fLInqykSL5MlO4XWrRG99Pe7LhCcQUm8lyatn6TBdA3AH5ktUOMo
iv51Mg8xE6Ovil/O1tlUzoLnnvsRNJZ72dvI9bSjK6wdVeQZ6UDg3GdERqnfkjTfelgHNS0LQFHt
C+m5b4uQ/28owhcizcqJooxqL1RjxdQ5yXJgQNdXFnkZ49Wkn4xUlHjdDsSo3vIlro5b5B9o71PI
/m79R/ium5PCdDkQyb6p+D+wnIHL2HSpL/6vnX5zUcTSH14B4SZ9I4PsicWOYhbbNbL1ESlw7Xe1
/Hzoz+H+I5z6WzEYsuU4cZy64LMN4ROoiuR7zFOj0Er17fCgmWJnx2q2FrEDKQQysKrUDl83ynI0
2ujSQUMV5h94HR65GPpodWZhmFJUYGX75OtgEteJX/bDxavVsDT3WpBl0zIOAKLM9zL/R04rYVGr
J2Ph4fm/9OOMNulSUNxY4siWoW4nyiv5NS3q4GtSWZv3evmq+BtBrraXp/UTMXZGMWPsPRtqS/Ff
KkgUZxabqOIUF954EbTI0avNH/gJVWmfyOiSuJdvFU9dPR0RRKm8YUqMgvnirSfNeJNWX2FyO50H
FgDDHpIPjSLs76hxngDiUw4QMdF1f4hysMLBb0r/Ipi+ykC8Dp0t76AHlnzqy4eW29DNMWy0PQFP
iAdtA9WrOX1GcXoTKAygjvseDlA1OKY4xtaWaMEdy1eaIfQ5iqQRybn+ZTPoK6suKaW+XQx5rph5
ZGVh1EZoVnLqL4UcMQdzmJsTUUrNFEvZJlZ/yL6fTt4pEwHtdcGXnKTAekpu0hLqPJWqibx0+AYW
m6iyW3N5L9UPrqey5dggxC+wd+O58RMBE8KzD+rMdHH13Ky0QdfWshkRu4hzFDFcFu1/Fknx6FOB
HbES41q3Yp7B6wufQXbQ4MSh7tafPq918U0xTBZAbcpfsQdKxSq8/XUt7Ypm5S0D0l2po+hCSBSW
BOfbrPQB8uN9HzXY++dOoEnS0jqQ2JSHB8MwdH1xTQJOp8v8jkW9kWzIiUpLoQD/mMEu5IGtiREb
2lAJ8PhNPyyDBR0sm/2oWyClZWDksb3a50bKh1aypaO6epOZ4jYXuqThwb6uX32YlKwE5iCHFAoU
tUDnYHS67dEY7EFH1oLSvleh4A+7Kr4K4plBgxMeRukr/Z0fUCCCWzUuFuk8HtQ52Q1mYF9lqbYJ
0JF00pnekJ4UImKdd5ONM6Q9AO6WgsH7D2Ii/tSZyG8vucKPYC8lb7Yj0uWde7jHoP/yHMMpGAC5
fGOoGTVguPVNGYQ5BVOY+RxFNzZRpgthRI1ApO1J//wZAZoJJGOz8bd5ctsug/Ypd55SZkyAPxp8
alzPlS2B6h0SrydFiLLjDCpPrRdZXD3i/pq75P7B6fzGxDzMb0JMQdeAiJzr177xguQPS2x+ISOD
MRNQXtcVH9Q2Xsr0hyeFcCpktsb4p67ScMYi/3/VEBDNt1Blpt5nl1yd//Xf0Qj+S7qVzLqgKKJG
28b+hQ5aY9a7/AmYSEvzm9VPFutF/TmIdNre4t9TPdxVvuFmRAghDreUcAku3KbPSfqlu6VM3ZYX
XYnLXoJXhHfjR4vMiFPOTjepDGdPml/hZMCkM3lIYbi8HKIBXwmcdeIiDF253AYS/fsxrC0f3XNv
/SPhHzMGh3fqvne/Oyw/Wz/I7/RMLft1b7qllN9Ui5k6s9ZgTtenqvH8p+D/pc6xCkMArBM/9yCY
5Xn1QwF78HLTV8zazMRzebTFaOd9tgN6krSMsNqjqE/8eaXN5hWc30taE2E/0ONzwoJ553gqwj/X
Yh4BRn7IxUcvpheeIEbQ/BIvo1oRIOa4D/ejtdBpmVDNuMQJ5Tcom6zg9b3NI3pAuUL10w6NlF4B
mXwbxtgLmJmvKidDijXPWqsR6WkD9PMNhm/Z6lmtCwFnVrqzN+Eu95yVmCHHHV8e7vz4eowXAt1q
MZmzQbJM0eulo6JZvMsY8RhNAHOlkam991U+fq48UzPW4VGskCb/k6f4cGAVAakZE+GEK3vnWv46
WmB9ovDnkhPGIsvUuAFzfHwr+pJZgKMwCr85Sw2e32HPAxOPAc9d6lu+PvF57jDSxszcIEFhu35e
FleFGkBeGGP2d4lQtfbV0d1K3GscbSab3kMEiOEuroto35UFVoad0YjWVjy/exqOmMjGKZg5hGTK
07VWmTIUtWD7ydDy3OgUgFmL/PEhwRl+8L9ucKGx+QaOtxCbLGSfpRQQyV4WPTjv6ltDml3RjkCD
CTM409gsMv3Xb98zixiJk89pjq935G4kgn18F23O8dUixvg574WHNUJasgrq9oYgxq2lsc25bp1I
URqXixu6y1wwSu3ms09KuDON0epGjXLq460TfCn0FSvDc8VpIf69F+XCvx33CgDttGhHkZJ7UXaJ
RGadGJYQDuxry/Gsyplbp3BD/UpP29pXxOpSO9J1gcHU376NLlH5tvZRv7xUnIO6Hx3U7FJOADT1
d/LdE1meGDj3z1HmkOf95pTjubckWY220cfCkC3a0GZtFgal2HtpS8F6oe0rwDpMokspaaWPUDEV
sjo+1gmjlSl6cwOSVkFU5Km7Lb/zwy9QgsjtDq5UABAZOe+0u5e8+CZ6inRRg7nB8iyR3FqYfn45
9SOrMKFlL2waBtv1G+ytqBSRXYtfGP/fNuK6u5YyJbiUYgTLADNzaZ0FvlKL4jDLfPYSH5CH288i
AKoWouqHWySFJpUp9ClUI+7SHTu+D72oE8JKaiC0dut0KvyHIxWr2NnCs0eWSpG9yBiXyQwIZ7Rv
UwCJ9xbGcrZuM5s9NlWYYWQKPnnX0e6O3cEaIu2j0ygyv5Q24nlmLTHqMzNlmm6039zeUIhVpsoc
FQ948Swtv0BJeT5A5Vpl8oT8cnpYjDi4w8/8WRo3+zpG/LiO2buGinxKecWH/bhhl7zRKOgGMg2m
jrLS9DNWZq+3Cro2SFaC94XAJ68Bi0phuRvX3n1ujsVuO0x2aLfvc9c1jD0C8Leor86EGLlY9Qxy
mL+dDAftSlFIf1FpLlfY9ewf0A9Y9t8L2a/Iyk9Av8te/HZDPIrEz7phRH6Mrq/WyuUa4wK19JR+
cJGvhdWSQJxiR7mqL0Nd+xs6Hu+OSZYWAVF9zREBpP1TZ8a1WjfI4TrE1Wy+WXOVQfwdi11G4k32
NJDwbzpxV7l/8vfSb7hDhbidhMoOmaqkf4Z501Rm8EDNUXZNpLsTLMVFgJj3Q7BRwWAf/hV/u2t9
a8O5NCza0ciBDR9oEIu3+F4omTBYKiGYMEqnZTJzttN9CAZ8pwMR4snbFc0m5ig4IGoejUqLbR31
hSYk4LOAffybdsjwBmUlV/NWWxx/hBHjk1uAzLsyoEyDVZKs+bkrgw45CH8VxFdr8efNashBvcnV
9WSwkIcyP31i+4fgp58gqIFpsIQ9Nyfej+UVOb7wk02eeGm6The4P5xqzki0YbvKcZi2bo2v2nw1
OqP6vpqx9BFgYNU/ZEsYNb3yqVi1icJBAo7KR8v4TxBxGub36zO0TyMONn7leFyivQem2wNaRbvS
0TqDYlds2N1CJhJeagjy7DTkf4jezClsxHwI6SQECcR0kS7tLMT2O4DPwsKzyOR+zRxN3lm+CweS
K5At1Jv08bKezZjjFFfOINYZOSt4RpFFYsSDrakF89WHhiaeeWkWFwv/kk6e1pvNzfS1jRYAJr3H
Aqz9Oz5xr9ZwIiTnu1U/vTiYfLNcM1PDppLSho4EtZ+pt3R96f7p0DOJj3hwPcZcCEtH2OL2162o
KaoW7ONskm0zZE7685/Y+F/cXzZSLkgqsAzh/LY9dAw+K6JuYp68HE4emFuQUZHfhUIB2xnsln8b
frmmaXjbHILmD2KHoYVuv0/e9sCfuAXn7Di+kv06WlP0kwFARltaNgSus4tDavhMNCckCvZYP25L
Qd9G//mlEHy+9OXyOhg3MkJOgK2n8kVbwBP4/pUWrbhZTG0qs+TpKzpQyQCGQ6fKeNTl4fPLf4nn
ZClSLDAaG+DG7OtCduiJ6kaMqoFmExeafW6YBlo4Dj3Hc/8u8yfxfKzkQMbQadlsk7hTdexUZ3W0
xNu5uOM+UVjN8AfQixs6k4bwbMbNSPY+P4GW2zAXI+euReY+zFBss2ITG/0cR0WHtLSd8Ey9V1O6
7JQ2U0QSX/yzHnMKBbMzIHsXt/fHuJCFhAmLi3ASETW4DyI42wpYz7WW+1mtA0gkKqeh2lKnfDUn
6xH/MHu5C6BSbeJ9xpAkGI2gz5p8nh8CrsV/wlcpHtZ8VMIRA5gh3d71tZ45deOJ9a9MXIrkg4YQ
M4rcKzFrRzzSyMuTynACWqRbjzqUuF0vDJsSZk2tCl8SWs2zzo1pmjxwT4n4g/u9LA8NFMlzJiNx
Nl+kTchUhTxDfnmcdBuzZzyPGlpLmxpbgtQuaAY1xdJDaqybB9dbbD60n2/h2njakFJ3KWFhElRX
jaePps6Bdtl2M65YeQRmq0lTpPKTDnKk2pb3H2mrr9kQLY6Z1tAjBYo2jxSBmUwBz6qm3pEbYHNb
FNxJCuJc3nUZI5Q4FJ3zBWLwnxPT5ZNpM6MY0NlIrhE2A+BS3Cdgv4HV26caU7d9VP0MbifitNQ8
UfpqhWPFECtuE4AvwWq6jepdROj3Plt4fAtZPJovweAHSAYZlBOjbTnM3HvNDpOBJ6NtMM6dExzh
R0ZCp83Asqnr7BezCeREBpD2rfKs0CMvwADadkdtWvyzgZ6IyMHCjtKNHWyr455GViVbGKjI86xG
wfc3Apw6KkbbxL8zO3Vi6Tk7g0EF/wGiZtcZoWSE2mnvCjdlvuWEgiLc/N1CYh11D/H0gSU7YSNN
UZC7rclEpPrWODIyZc9VW5q477Cw42AIYoK97ZYTFjFbTJCObULnYlqmlXgcdIRPV82zC3bdK287
09/55jXy9ijUsjfWryyzAgfpG7h1xxLFI3LPtPq5AvjphsGkNrgdPAuYDdp/y2KG/NrPMLu9eey1
44X0huTuO2SDrt1yQDdAIRcve4qCQ50ybCtWeD2dV/Pgyr67ZNtoV+cnUHVFOXDNxF/BuEW+VGIa
6wckLjz5tbRmDm9X8eLS8ITemEokbxyZk0wr5Fol8qNlLF10Xc9bGwZZT2IXKKPEYybWE6F5fXC9
yS7bhVit/sE3B6SgRMC2DhHr0tDpYcCfcnaG23yfDeLVv8Uu/x2xf6kLxaJe8R+aOZcBfSglvZho
CPDKmqVGc4og5VVgJv7mK/S95BwWDmeXVFbHtYzZitQBucAXSWawLadU1wYuNltkM13raxdvWT/W
y7Nl0i4E2MoonrSdDRuhDQ4WT4yOTS8v6Nbzi2GJ1z2FYTb8p1LQeZHJW7EXrhMgeP2fAJ+J8E2V
5YWaF02JgZNqsNKYcOZq9KW872Kj7km3Oo34E8K9Q9IU6SQspSZC4E2JHnCzf0iwEI7vUFroeLLI
zoXwKpKs1UvGM+jZ1gG95ydH7nl6SMyD15KaINQ0Y759LyqBaN/suPUnuKj2KiI0z6vEOXQaC1RB
ZklrljTfjQnuhqNrWZiiyMLZIX0+WOOtB16ZseccFgvMfM4DNF1TfqIojt3t5iCJVB103VoOYZ1+
+Tose/fpQ78JXgLJt5YDdKJX821hiswqmcK9a7v2YSomwh5GT8/ErPIX73q2rFEOV5iFclaY6NhC
W2MQsBVcyOqn2qjCqMI+zlN4APcultbHk/IVQLrSyXl+8PsjnhCsViMnkRDUN4gvMaXC681LhX9h
GdSGRZHs2MMJKgDS+rAyVhPlziBhR6fVkAnyltGLUFtfQyflMUuUD7EtjLzByWyAuYE+37bsRQHU
vYWPSF/eKMQOXuEWkgJPlIU9j9VSglBqDiKtkEijcCP4MXuMLZb/4Lay4u5dTnwrw0jNMgY5DU4h
BTu7xNDvghgYQNgy729ro/dnGXTk4dBWA90/FG4ATG6x/IGQtV1QsmFY7KA1PY1WTyotlOPsILgr
z5v4a1PlyZjurmgdV2g1yGw+J/MOPuxWCEs0JLpRjdijXoB1CLGgrCw3GYWoTjwtuMtLBO0lYs9j
V0JvI4rCWnDT/D4E6AlUxtIjAFqkNDNdqt4vTbWwx9APKL+f2XenqC0wTHujSgHnkSwQUSxQ0GeN
3gmPWZNms76knRh6o13usoqHoveM9zVXUGGNnBplgPgrlR+5Ijn2VSN3jsIeHQcao9XYv4sEMsFO
UghPsAVJrvhX6AHRZuTYLeSHGhPk4YkOuQSexSbTF5W+YRLqA2CW8ZlQDF0RyGTFq4g9VjHySg2f
pC4mmS98iimn/OHMVD5EPUqy9Mdc2bdaNA3rK9RR62e5zo0JjefdzXNHwM8UP+4NXyLsvPqJBdC+
3giMkRipygL4Fiok12HN23rM+T3mhnVpYny9KBauMWIIbgsG/BRkOy7JXBTNwNNGNi/TG3R7O8Kr
HPtIb6a5bCSKJmsbDJM38w2/YQdqSGNmpf4zPo7ESSQtia+mnbyznMeLMtCA676SxWuhRYP9fW1g
J+EOR7NhEd5euJ9E52AZQtChSTLU3Jj6t5jLx/LN3bMcmwuy4WQPSMzCzPQ4BzQLXZz3K5svVD57
F3GH/M2NeFALxfSNuWGYHaFSdPah528DtuFlS5+b1+gg9jkuHX3hhpXndtLYFHOBW8Y3PF7fjFzo
dYZqqcIhP1XVuYnYmG2lLF6srt6L5/CwcY3QW5NyzceUb+5W+DjTH9mQlMh7OOkTIz6ulgPewo8J
6mep824CmwF5OSbZNQH8RkMUVTKD5lVO6/UJcVosVjNGm4002hRgWs/a7f61+4uB3QICp4MHjKPm
mpVa+Q8Wr347PP00slNQN4VCm/6OSaRZ1+BlbdgoEKDXcDW4IAVzJqsfa4cGxZK0jIwzBxQWG+p+
BoFdm+jWGtCyf85c4w0S8dGNgTE0PHKFx2OWQX4G1/NkqJynqARriSvEhlVD+Wft3+DBDn7Iz5nr
pUtG56N4/qoOCC1+od/3MopO/y4Ud5WQBiOgviPQ+hBGaun1GiM0XtZKz2c0Oay8hR4KvFetdhsX
qgNfnqTaFyl/ssCLPc/VyXyDsWATsiDBKtfizLmr2ICANzGUQfoKKvOhdjHB1nSrY8fgfl9IwEgK
aTHWFnWI4iCDriVq8ffp8sqC+oDEa7rNXj+Uzo85FFKkZy+i07/6rS+VcV5QXQ3X4wjO8IPN6CSO
B9nTP9TFJneIxZ/90p0yBSpCem3miSwTDVTzgcpQF5nmBPyL9M/dQzEYQR3tjHx2/agL9HRoXj//
pzvK5kBKE8D8noiM05Ce4Fd0FPX+v/NMU3oRAb0Vw4OxDyNb3Nl1hMIgRq3cZwKN7kcLD2Z33slz
gFOYRg0XcKW9jOqcKTjTtscLb20LWQXGDtsI6AhWVssqMdvbgE1J0P8ugOS95B4zimDUPJr5noBN
Qe9f3G/tv4ESieCaHS1ZInOOiVf2UQmfk0DzsLrVg3188/IvqSoSMBZt7DsrHQG9ZSHdj8hXTg1n
ujj1AbcqXnQguBuDU3aVfifUjh++pmVir8XOeO6VSbIyGWplUl2hSHsfPsrslIELIY0YGG1Xxv0g
tQekJkoZLIvg6nekxxOiopEUScKEe8mPduPuL5UiVyhDb0ZGh0CATZxKofkgwkqkNZz5TLStO3Gr
glzprjfyTSzsKaNne4ZDYerJHC9k2SEWWY8PN5o02v/7mt0DyhyjcKCQQZXP2VS8Bz8kHzishRmz
n1REANGEV+9T3sKh9MqWsp2eFCYlKYtFjp9zvWiOLzsJ31MWAlIQjWkFD7AR2UpL/+uIJl+sCyJ2
nyWRf6G83uF41GDD5K7DigpAFgdbktx5cygCJbp86PJykyrjwjWIId5N9nJ+ZAgEkfweIc5vjoV1
rctgKHfow74xvfWK9LvGUqmHe9qS8Fled5Cp7HXU5wPgivMCF0lgnhjfE2Ttkk7/OSAVsEE4Rvhz
S5MEBR+R8WzXETMFS+KINV6diOpW1SVjcnNsdkA3GLls705u7IYxsBiGsUCz4f4LXM9vczWIkau0
/ObIeTBwO2FXVOV0cncxmx335HrtK82hlabnalKBKajf9z4Tp6N67iRbggAi7yv2mJrB+QSfUfaA
5j/PEmk9UpQ05LRFXj7IU5agK9GFTBk8bRnyNJTcOzvTo12aMWGjeMT55CRdQ2B/nRfu3SWOzZsq
/j9AV9HmXTYtoFGh/1GmkgAuhYlWDR1D5Gv13F0KTN7fXqvV4khqcFIb7xacu7c/spe+pTwFSo9Y
GcCZfbJ6/ge7FTcaD0TsuDn2j/fkNmKkaONcTlWL3fuiBEqNsShSRw39bkuynIGbPEeNXzh6Dn99
NYAnKyodEsyZMPHhYUAH3UIQLmzzDh9fDmPjb59fR4I7OoYcB43tq5N94wwST1NQV+/uUogYbJN9
7q8DgrRnyewXSdshGKke3Dadp4dMUzgZ8Szo/jpRBQck6YnQm09XFwYbK/jje6p0QabQcJpO2k3p
cFGxWcilt7SjaYe6/FQu9hlta/NsXdMM+FJjwJBrDyxyKr2fNkGgOgXqr1vfOtuSK2rSocpTO76Y
07O62sNA3/2C5srAWwRWkHwkTUbO1njML+imMYUkElkw7GrqGmutytJqb6cdRT28bbdATIkHiWKt
VMEUr3GvqMF/b5UOZifAz48Y2GIuGhYJK8CQ3cHZogLVjyt6h1DxIvvR5G5gv/3PSUOWLqtbxckr
ObWTi56d1OkgBwuyASpoBmlpNhBH3Lf6FhgrS/UUnwSqy0y6o/89y3rMFKIFOwFNVpRG7YXuCVHc
k3z8dDzXsZ03KtFht6OvslD5wVIMU1RVtXMMaTxZk/Q13mjXHIQC4UkaBejT+/qidje5DQMgyE08
8Q4DTXwPYBydXKz3NwP/NDIg2v/gGHKL3FhI92dsYEqNPbgftvBJP+bC1VIXM8vM7kGsr5EcqaRt
sAc/wQ0kNQn272zBFtaS0crC49qZX270UUpZGXmRJHNJfd1ZeQjabodosxsmBzaXxLTdLhWurTmy
FSgjHRF9E2vy/bppBB8m0wbDLQUBTCuP6G+20yKOur31ck6/Xrn2d58Xj1leceK3BRO/nywW28c4
ATMcCzaPtDOatt4UnhgAezjc5dKcdQDE8UM2/zC/TMca26thQ/4YYPGhrAqzJnGuldTAzZVPQQIp
4UmOLu2eRBhaUN6o1AQKlCerehDA3AXdMiNORmnvcEMt2ZhiaI3JuEcijVEYZWlQE0NnLBAcbxT9
yAFmx7RgElwH2zT3T9ew6LHImyrF+XnZasxvhp3NXNu+qeRqIL11wR8FnKE1i6mNLNdJ3SHTDHcg
n++PuIW0MxiMLG1tzKI/XKp6JxHlDaoUL5chuN/Z5PIUqqyGgAfPxsieFw4toUofNM48+DZVeOlZ
OcKLGlAZtqXqDgsDfpdziz/hz1oLKyTC+LlIunKqF3cW1G5UBbCdrFQa+Gb83acMHptdj/RtKpE/
U8IyOadgb5V/XwBgWszooLq4YJIuIat61PxXCqBeVgCsjaceK0oSRdY4thUK0n4Q04YFfc5C3mTE
wuVfmfb5A58UBzQomQdRaxka2E8eKAktCWOPiy0b2jU5zl/oCuNUvjJIC1YUN0AQYS1+0jpr2R5A
ED5jkz+Nb70hJnR6B03hqcNrTWy2baaVSO1o6pvhri7oLSZjNQUHJ9ZNPS3o7SiGOg+B26YL+9nu
ilhLaU268W3X3UtEeiclzmRn1Fm/5hlBKOyGrSprSR7rD/4WOBgYhArpqV6A5Ef4+/F3X+6VQyAq
EWczX85Ae26Tealh8gTYIQ1qtY+h0PNOmIASHJiRdJt2cSi4UAHBn99IgeBOk7lukrrKvH6iskwX
hHTtVmOAqFv73+I6XoNLQIshb1BiZ+yWXdjMTgzq8zZuYhWzG8h8hV45R/zWBSnsX339W4jiUdm0
bvbhVbP0cMJ4lhEhX3trUJhrWcsgfamMq3v2a9GlGQOkyuxhG68E+JL6cWuKlRL3j/Stj4NUgh0M
DH5yehqR9hgKA6qIv8MLb5zjBPx9rzqIn1pgArDMa1Rfl9ErHRLZiejcVWVzyP3rv8/lhqta4W4W
HRZh/Q0gPg3FNhvNaVZe1bzgTqbmqCmAnx5p6PUNhiZM3iFYLCmyav9QNF/ebkHIQY7ASztQ6rmS
e/nitNeJL+svswC6GPKCUdsKKD8raKOT5E8e8/+6f8AZdSNfUgEgJh4iQaplqVUHO3Qu5BuRh8tQ
sLqZwLFwaexvbSzeC3J+YbqsbEOszmU56lhnppyDlz90pJaZFLJK2vDqQBl6oP+q0It/zeG8GY8u
znX5ZsDFPX0yurNTtv8JEW/xVqu6P8JSxkGpwo3lhXCWcl2qFla0EPPqK/X8/rKItoYPBGyXtk1f
PQMQWRT8YJUlMBwzq/ahuUExJt79p2+mr+EQtnNpeTc3/KZ484in8wrOyx5Q/0ouZdRlcLwwFtLu
GpmUzbYsKqglwoHFlsC7ZUxI8YFTuLJRV55k+RTTMvmG5ToMVplKbIOGwU+6KSFADRIt92bhBRvS
52ksL2i6zl2+eTHJam69uNP0Lt5LtTfydu9TUlQ9UC5AIGZ6fSihnexpV14dUl6QtG+f+XtWUfys
O5Ha8qb2MCrKRx/0EZxlivI7NnqD/YBsOu74NfINMdV5yFauZJf1qTwyoOGRCS3d6it3ZiTvkNPP
QArO2kidKDV6heUHVyqte1/O5bdUwxkHmzSU3HN96uvmVS9xhWwIs/F+QKci7znfBaGTy2yT6ktq
W30+fgdh1AuHyJSVpu8HC7enCEJN0jD4WeC259+/vPhAyOv8FHafAVvRWkskPchbj/AYVRBTpw2e
x585+IMqvZTq3q0VuOSOVnit2nnDBCrCIk+ipoxGO5EWjZ+oTJVsYf2Cahl+XNsAKbzGfjDgGKUB
QnYKeOSueqdWPaAVui306HvAL7QkGt85AFl7O0PyEewHhZLJ21SY3IZL91PflOzLKG6Dryl7OKzE
mosYmW6wD9qazIvkpHRggT1dq2ltvn+dodBKZdxEjiMTfB9nd0yTCgjBm3ydtssi0iJL+Y/LIImk
rW8ttZlgz2MmGitYJYjI6IoY4A8aLV132qDWBNWtDTTEbUHR8R7HovVvIzCvPlhiz8PxfPeH5RyT
5vqc30iSc+igsmGhA1kUAPeLfJaS8msDI8u/tU4LtMIGVuVvucYRr10x8Oy0o1Vl8pt8taxygnbh
KbbAL9+vTzwkgiT7bDdDJR9jLKpuA06vAS/waBILF46Tzv2WTHYzpZV1Uo8n0X8UqPuTjXJIg7b6
knypQpT/eaq4R6iPhdRqy0SfqLZdGWjTNkzpV31FK5iKEbiYGf01hLWkZy6FZxLBQGdxb5d4IQS1
VnIdAiI1LDlB3W2bgWq+6ltvlEwbxfczG2nHLAaW1F+L11Sz+4Z/95NlXuQPKG1m+ULoAcHCPbEm
XVCz3d69vogoF85k75D91qbmhuTgm5ShKCWb1fdla8VBIthTKGpkp8NAvQFY6jly3cf52zYPRO18
TOHHCZOw3/aiBb3AJSri6OJOQvQwm9trfVhKNT3tfWKAiPbEKXhtuG32ooJcqxNSWGkJSg5EPlp8
JMuhr8s+Hx74IK3X0X/mtcNHAAl5HvzTOEJw51DZ2Q77O2Nkm3wdONjWxJ+Lloq4pKHZK2Bya90S
Bf/hyHkuaUsFWJnUY27fUfaJrm32bdmX3Q6SLHDgF8fidDz2zovtcPorKn+Ts7a/B/oAc9KvQPLW
0Goj7zLCH7DWtjy8MefUBqFhVtn+hlNt5ZQyP45eXio91+pPRl/Zu+wim/JqZDjacHxcrCrFmWxW
JJLtS9pk/wQOenJ+qdo1LvzXcrxKePYhuB85Cu923q2tcaGDHPVCWxgADL1khWKiVnSZtK47FBOe
pRntfQUle+NB0VtHFKGQ3RelGlz8FNgnsE1qBFk8U5wKJ2XgEOPe/0UvFFVhDfRgI9Qr5gn9u9mG
m6aAynDmaFrjfEa1+VpbYk7DGJZyKCtdBU1Cd3F3IYDfUJJT+VxGszAFQ9QS+fHJ1qkyust4cZ9m
NUXJPwkxFdNce0MPaftoRffkvUVYRdU3ULOQ8mlNtBgM+rCVnzdN8wWfXqbkghzsUwpVzo3075gT
mmx7i0AyCP3J1VBl/LPPm9uCQPWd5iWtP32Bh1DVxtniRxAGDyx7pmQfP3lIMDGSaCxwzWk+T3QN
UydmA+KHKw3blikY8cDF0BHsj882ItQfgcwr3q07h+TY8baTKQmvwkmyUKcrDQPhGy063cJYv+tx
5CTbShOl1HEYj9oX1wW8Xl0wfwozThRgMoFzCdvZjOYXFMnJq7mNcHnuj7Wz3vCpG/QEgpKbZFa6
86m1oDgAH0yDbTGnZM88NPOLxVTtejvmmkn+XJzHr7sn4cyrvhp+kMfZRhp9mxTRppMZTrGeHWc8
idtlubF9SE64m+n7hMe8UdMwt7x+QSG2u6qdeNPSBiXBddLMTlpetev/lYJ661zSvAN85PeQCewz
sxz2d6r7wza6ozgqmiO21d4eVTdbMTQOWq+otVbj0YN+fZORce7/KRtw1ufw5OAnZHDh5J/D+IOc
ff8x2V9hW6FAAT76MDijL3vXXiF/aIQrvYrY8Ah+yrrjLvWRBOzEisv/0h03DX/BpDY+1fuGwEJA
eu3MAYZcs0slO7Spv9fVq/3G9sDsHQYx3iTxx/yFNGJYdsOCTZOpuF50fmfzSPg3KDyTqTuX+CdG
Mt5ZJ9/z6TlcU6fMubM3nZUDbLH0EGo3rk9MYmisgl0FihKLaOSYRXnzmbfO4tCfymTJ9s04oRwP
/zRjutKsovCSqEKE42tORbzG6fNKh+AgERWPRPo5IbSSPwm0qdUFwkEyBKfjbLuAsclqkodwvRGi
sxmbCc9uwPLP+rmv6gP835s6LJmPgePMxL3vFimbBqGZ2QxOcPXbmpfpOhXOv4IVjF4zhDsvVKj1
oZmloYjobYs+IpiRfl7F4rLFbtnWr05jayt4Bl4dHbvHT+W+MoxXIS/B75bTADlsvJRDBdMtV2+Z
B6KSG2aFqTb/YunDOhWIwEiSsbPWRUSildoawKDGbyhPbHWMMVpUcE5cwAWTsSJg1FALWZIWPG8a
I7z+ff8BFQhPu0B9j42Do7T6pF4Bwexbt7nA6eivcu9xYIFKIMR/jIUhWAW+mgZLU5gMf6Q2N5xz
StF23x431IPGcdC+yVAOZrWvpDN7xLTGnAN67maZz6uPJSQGyoGbaQ2iw3lYW9PkawLr47u+KLib
fQNAbgJhAQiacexieLACONFwiIAaQ9vP7wEBQU6NsBsrqWwXUY92Y5bhBn1wEub2I0mwNOICr6+m
EcpiGFbtlW9K1EqOn54R5kRKN/2eHjRqz1iNRJLOES1TVeGq7QtTj+O1LgmYqgVs/Qzg+ShoU7UG
zRSFh476q6FtH2nLRJ8OQW7R0X76ia7EW3qbCaeKChUA8bD/u+D2wfgRKUUh45+FIJpD78kmYKxk
rwP2RWe9c3QNVwnQUWAmSp0R9tp0VdxRHRXC3IMBRqdryyA+dsR9WDbjZZ+vGvD6LffjippArfhF
7ZUt6dCKRQjIu8rHG9P2GNnyfK3QK9hOV9MfiC1KcPdejtTPSSUDSudjH7eNxKo63Xk+uZOgOlet
orssHi7g3o0YcJhU511DX9nI7T19l26Amf1ECe01ioX+S43SwnK8YBDo4x0IJvwM9vxDD4mv/Cn8
KBrmWKDavn3k7slsv+rcRD9T49VQ2abriLmkDqB89WOQwTgCAjgsY2HooBxNaO9aIA9I3dERnjJ9
Xa8A2wfOs6YJN3AwwxwVnimTfgVHspjCVhsEdbczAv+9DGEwSyVW9isNVW6brQJLrti1gHVLxG+B
J7jBWniWsCQqivOoVIYDfJ5h2/AhB4BJ+kGXsKhwOuLqiH+m6L86fgbLQkzvoA0UvF/t4iAeiQ5j
bMDM5+d6PcYvf46nf6IzIsQ2p4hCSI94x5u+d1E3ZN4TOv3+oKs3xRJxNLnofhhJLvfZMzfaOFJt
FpgJ7TyV3mr58HKF1KvjwyD0SaibUDTxdey4UTGneX2m73rDKOkLoKoDuVsOWSO48MLanL57NP/6
PrbTqaQZn/TwErOPgrDpUhjyAtxZNSXQEnkiMpJ3wn/Q29MCtFSJVJ0LUbBpKKnHKJEI9mYqcySH
8b4Zgq2Nlv1Xu7aRTE8oN4bGQa3JYfMFTCz+CSA5QciahtIVhPlgm1cwVUlHj1ilyw8goKWvMSq3
/h/yJxPkSXhO3SW6CY2UN3NtioHPuYWO5y/J7YYvn91aGIaVfvnFrxmBUeT+4uFadG9bEQ3tpmrH
iE9YvZmRtdwA+XIrgIvfcvfOzBgLtIdKG887nX/UXYyshfGzprvsrFeghZI=
`protect end_protected
