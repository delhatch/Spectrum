-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NDz3J4TGuzpBUilFkfZcf/Z3VKZPaaU7l3YaGHTApVM2zT75RV0w/hk+YDR+44z2usXklfS88Xri
Dux7FW2+tqS4ql/QdMgVnP+PwVuF6EgjXhnYKfLCqzsLaKq+AGc1LQQSdV0h+4wlC9u0YNWd7gAL
LSsUJNtZAoxHaV+g6ixw5cxasfS9dzevnoecshIbJu9J4SLrs983emnYqhpgOQatsqxvAqlUSBXX
WeIeWK3dQeJSqnlWvPeQaQEJMShac3+yviZ/L8981EJU6rVQ3daiSBynUxrD4kQxetzXn7t/vOjI
4+xrUrMUiNKdMtFxk1I+/ljcEBQiNCh0gq0f3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
lDJe4qleFcyK20T9sfvvHvobR4GyOVAGfDa1YbHt6Vp2zIdOEr719ZdVymt1VvAskU5X0LsA8YVJ
6wGnMGu7Gl2sAdjZaMUW8wXMfmwsaZS7awDbY5MXnA9YK7FpzL35PMbCsQrnPMeLA1TVplh5cXQM
DPkWqjm2jMyb+U8tFiJf+b4DG5LywDwpFRxJ3eDAvzkoSXEWwMApD7lqjuGwDadvbj/EOY1sx7it
viAaK4BQjyxp+Noq77Fay7MVpEtx0b+iagsNpZ0gQaOYXy2I+ZfQKv8p45DxNKU+99EMREFVG9Y5
RpptcH+XuyhAvkbv4fhy8baASRBjRM9CUVwjDpPBulmcV7OwA8i8lnZ3VSFx4F8h4/ocmAiMu/92
B1VUVyejStvhTV9NOevCtHbfEXMEceWX7mdoU0/oLY7JCMZn3918E/EsJf9b3DiOvG8mjDakoaZu
+FwZKTEBaKlQGpHcdByYCfTqEtz6zE28yPiigpr74Z8OgvuhhIMVOiPoD7BsQlV9g1V//XO5EnCM
VGHnU94f/ySBFOy7awVqi4DrKY8134tA2J+aznQvA6CfFAJRBbMcsTYqZEJU6SdnXz849IHka7Hf
6D1RSJYNzGg7xCreyoLjw1mtTRqFW/cw/x5PhR60mseu57K7vffsnbzJWqxgrBLUyGMRw+S+yDpI
nu86dmSefcJc5/SrPi4C/1gfXbNrMlCze7wtCZdnXxAlVEYtAHm4te0WqXuRfQd6+ha8+eHdctRs
jpR/vtFUTiG5WnlHHccwZbMpSiyU6ffjb6FQeov+a/2g2UoL+jWFogK1z1f718atuqKHaQ6notaU
2XNHVKulFJSthSWMEYSJfyyq5JlMXQv4cZrI5XMgEVwfy0Taj2IjQiMZczUVYtTKVpofTPH90a4V
B6LCq0cD2mJsdtqXglMg5sL8BUFPj99jOR16uSaFwGs7CZjuY/X4OmYzAPRGzkIwBNruJtKWeX9g
XX6nbREu30fT3b9Ilsaf2K5js0v5/20YoayZj3vNcUCMQvGlOdkCbOwbizYt4GOARdGMOhrUsNEs
5aVt++NJLP9TG+DcEOkEfIKctzFKbwdjm/uhiG6vd07fP9ZqSyt5IAWdde9kvHh2+YlHdfXABZek
5hZ7sUl32x6XRKC5FsLPnUm3khnZayLzcFeh6lnHV3UzWK4QYEgehFeG6Se6kqnMtoVFhS1mdpAM
VOfZIk779epNCdYqOC9iNQXYHuxROQQkU5fk8HZMHYDdFMItwjrMxSPiDOwmZtsLy6PF8EKiUmVU
Wtf3c5o3sz/nG/q2PHJ+2xHe6nCr1kysacBKaLxM9wXxqEGNV9AdNDCWP8LTKW7zWUZy/iVLZ246
POigPU/Ah005bnKWXfc+KjBrptVNNzqseXQI6C7665rOZ6c7d2BwcWefWtvHREIGH3jfjD7m1PZr
VqjdyhsCwhLnsfQCJaFx7saxu15ihWU3fPz1+17ZU7rMyQ8GpsxJygY8as61uabNACo+j3CXGVcn
luntGVGt8aG4mxUCzz47VJS5KGZ28+MbMvG2QhJfkwS7GkgYP4mB09IdK5Al5gejuMTIUkb3T5BT
7NwOEm2EuSpWqM93Y2ITYxbFYC0iVx1F/jZUDCfMfase8K65ApTGJeQaavd8AUOg+n3nYGCunjKA
NeHVJVd8ZhE7ITwsoOY0X0lVG8LRvymFV7PQE5B0Gktr4fb1QmvF4hWdksXypscE59kGoS6cTHWy
qia2lcReuquJihTBkuKZrvZZpKJum1AGgQUcmb14noWc+zHFaQDESlXDPWUyqCYU9p2aDAn0oBAH
yvX6YKgZSNpjwxb+8HeaOV0xccclWhX1pFpIq+BpYHU2kjz0+Zra81jxJb0SggUHWvEI6YDkdc8p
R6LRBrxH+pfuzITDoSKaBmimpHGx+6KKLfZsQfwelwGTEyqSEe5/YkxVijttZpIESGbt5IWX69uV
ldT2mxKSZL8h4NumVecnUrbYgaDuZoIm7+Fp9BbAIWmPrVkBhKoYR8KcZltuMGkY5XMp/Lk6g5d9
3wYSpbot3bSxPm/K9ahaRYdoMooAaAEFuXT1czh/bntcX4J0DOuEt9VUjbZOuB8AG/DYPgfV35Vb
UKMGV9Mw3RC/hr4YRGfOFACHphzhyCx67Z+5nZL1ZHlYuj44iwxWXpWa7lbZJfOzGz6MjxCqEok4
IalkbIpdvu2/TvfKS27nTXsRQgvSmupj79KKte/IZ7vbAoll4i1zHe+54Qr+9D625YBJhjAEhxgW
0Q/HVwYCuKGkyCOfJtO6v4uhFGe4eVi6Mt6PqzJsTABaOrEzPtI2FL2zB0Rrqt2XVmOF+KoKZF9u
bBHJ5Bn30YYscFOZxVQ021XHUjjSm1/SJ57oFFWdymLKXe7L/hMIT56ieFCLZx7UWJIQH0N/s1by
X4Z6lO9ENiv0I9JiUdpmYpGNxhSDk3h2g8b/AOfRzFoBQbsHNXWNTa7HuN6bngno7xIUPfMVSUOa
oYAa1kPaJe9sCgLGPNghaNPLJo1xPYkEkNtCjfJ8y+RQL/fDO2u6JYbkuBRrh3bBsTj1l5dgpqda
L909QaQ4WXTR8NoWkFfjQVUcjhlat3PrX+k+u3s9pVpgcUGA+quSPS4bOPfFrx4r9y5Mrhe1C7BR
OAaYbr7FtzOQdj2gRJKxPInI2PHKC2tJTpyhsfchhF2Bf9DXtozyz9KMYToF0cGJSNjiLTSdQHTT
lQK8uwZMbMNjk39bclRuuul3LR4s6JHFvHI5sPUmgJKazLMOW7/PsMYFxMLGUDb0GW01hgvCG4Fv
CRCrc1Sw4Rm3RX7/uVCXuHmWLwpsgIu9w9ss6o5bQ2OlPV2RQI+Rwo9coOWN2wqkqTeIRzqAlR/J
DTj1ZqhfX01hWiXwNxAEn0H9ZVTMTLSx0CFrCf++eCHs/YfCTEVBxKeePnfzv4m5jm6ah2X/39W/
M/GBFvVV2lSim/BY50YL0CrAhyVYn7ggfTGk7fi+gNahHYtUL5PUYUHx1+1kx65eOYJ1+cswmn7o
oOLFfUDSgCVk8cR6UID/hzdfTSBgu29B3/Ur/VLHGIfQSCa8T2dtIwGXuQQVG9S2nIwZBQ0jk2fY
xjjqW7dEIq2gI61SiBFDt74z8PHP1+WBQyiIDv3QVgSIwoWWeReznVuZwaPQGIZ2ECJ5Dth+O5OY
51L/EF5ZzorMm0QB09mdl/7n4nmkK7b70v94VVNCrXgZ4NSBIfC5Q/0TpIJ3zNOFP7R99BTUHEUY
CtgvVoqeCF2+sY2kwnqPVupnWxLF0uCX99t5uZeIN1yDss/+UMiuHQMfcCPyISugXvMdarzWTk+3
3EpTVCY48rPxbFPAjj3CyzNvVYv4uh5Gsp35wbjLKvWdFNT8Osk3dsdQx5sCtB5c+Z3/QxkC6sIe
0vKefsDx7i+M/zS8aQkCXHtlDcNCS4xRxKie7eN1ch6JpNCXZzeS9Gwj55v6LFCVqiJQSMe2lAwi
OjuMpjmogQhaYm/8Rfeq34oEYnGCo/1otCJISjUvL9pJ4W9IP5uxzYu7PnORxy7T/gu7+JY3wFNy
V+5EO2e3bbVxw5nnJrcPB+CmdQy6Eo27L2l6XPX6NSqcJ7BBuD+qKlZR2kXat2Cs7nCCQxPX145+
TnsdoLTV3avlR8UjyVFe7ryRm5l45DETtnZITJVJG3mkZXKZDiKe67bTseXknL//p4n0HqUvtRI+
9UgjrTBFpC+Zd3qWpsPDcdtrGL9vrlCAAwVq8+dP0mEfkCK2elez02JJ2jLbXP3DqvBZ0zA4TkAr
A3IKDmBX1Nn31hOGlHh5Vr2/tL9eMrw5FaCHn19OBaRMvlNPlOIhpF+Tha/l6QSFNLpeTcyxnLX7
L75MI4GWgTLmjEV3Y6aZl/dpGjc4V/JILSmx3WvVGvNx8xVOZrSy1dPQnu50nG0vcbTZO0aywv5T
TztVBpgIoCidJdhk+28ZgRaUsz61OUeQbq+EnMoPttWiXgSPB+WXQP2h5xIQbNaDHFC5JaPALhzY
uDiRCX8V7og8zTmqgIbV+4DAIE1ejgra2RTWg7xJm98cfUx3gXbacOb3bYluHf9AvP2ZGYoLCGMt
2FHpJgJnaXRJyPuyy65x5a6hhb9byAm4sRbejBJTKwYLUGDBGlzIA2tGiliv6EIdLw/i+7dNb/s5
+8/PlddmXz3VKv6Y6Vtlj2S/VXloB0U2aVmtVZPaL88aoOSAvNsqrXhmKXFG+Jl11T1Cxa600R4p
VEDUfzmxz4THQr94H2b3NMyHh3mFQrO//D4rMv/Yn5vyiFBXG2JDmbQRVvnSeT8y2TBl31DKwNC8
UB4bzhcOmO2W7zvhpOM5VYctdJ/R+2aVQLTq36TvST/agwmGt+GCndghrgMsxSVuVqZWLJi1zus1
LY/mY8SgID2anlrC6E1MxdDeSL3vmkTZN7Ez+3j28AFfCkY2wMhn6qzVpzwrv3QEB0aIzEwvaTS9
QtZxgajJFjn/je2rWxL6VGOTpKO4ldCAG7+1h+TEhVzOgBxA1nuzPoewViKIt5r8lkMri3YpJdpH
li0DoupGioCmxT5B8y4yQIL26AsudyDMDa+KdE/kIoo7Hg2dCMPonzm2HZ+4D5rK88vUUZjwW9TS
X45k8QYZWMzR+G6rDM+O+UMj9BvatHdAAA31sD91+2HsdFbTtnJ/8nA+QL/jNNgLk6YS/iV8OoeC
uwDJGHI834Jub0AFCH389a7Od7kvn+GlQ7OwU+773Vxugb5xvN7e6BULAxXZKMuGMBEfWHMx06sj
Sxdxcv4EWcAP1BuM5saVvvamjJcQb6qROOR5KmwaMkQPZOFO2FNNpcDItVILw8v0k6KXLN/NDurt
SEYARVBI/hVsPM/TNEoDGml/ae0oTt7GJ45rMZJ0JquWO9CYA/47LgvkuVxvpL6K8o5Lq5FKrF0V
DWJEtgRS5ME+uWd4ZOs2uNUzeaYO1GPjifjXY+cL0y02Zns3JokU0ji8xnApozU0cMR8g7b0oYkC
iW4zKwdNSFlNXXZNswS0UlTBSB0vqD5Kj3YaA/rmQbagciJ4QVc6MfWKJ1zOUBkxD6KyNLC9qSmk
Vkp+cCZJWQCyABODU3SY27+cM3kNb6GrR+K5DvXIDikNjldskffS7e+oddNVyMYXrY69kCvZgo+W
2uriRKHzVMNCB9Bx9XvJPmyU6zTEDrhCcqt5EiO2OXSY5fEyhz50g6Lsq+BDfMkhqaDOAuwaMk1/
jjKaPLHZjj8WV+ci2RHtadVEAyYun6bPjUZGh6d/i4eRQqbzHOs6qFlU7i/8GmCv6ey+jfAf7rLu
5LkXbc4zv+NrK7WtVGa9uLoVl0KyBJlLWca9o3eI+MMkcmNVjY6samijExhp6sEhMk3I1/j066Xy
ik1UHJe5Nv/pWAi13B19pOvM3WtkXFaZJnYTZtdtlUS62uFViY1lwNsl94UUmSn4h/R7PoVjmwC1
8Hu9y+ZP/Mn984i4wfWLlxWt1UPdy8nJmS3ahVM7ZwSBsgUYxufC7xJdE2W9jfWoftevTN6YKAAm
zadVXINBeZISblWz4bH4i4Yyfi9MwNrQWBDcH38DHfJRpFsuaLGlDQ/xRTYhQGgSW1h9sSoBgMN8
UFwqRwmlcAy09j9O9uvSHEjmh35178uQKJUKmsCpmjVGFzKEgHJoR6slJbmNl6+qNChTDCzjMZ18
dGOFOAzJk2xVIBp7RPkD7Yn5wtLYs4CK1Hg4HDD4rFNjBJywAfXRU5lYlI51b9rrNZcgADVCyBld
SAyRR1sudgkh0rRXG0QimwoHUuygle2qSNJXTrB6rb3mSIUI0K1e1jwnfkPslb5GNSHqocftDF6h
wF0QAFwcqEU7Mu+llWyH9IXJ7hASenL0XehvQQpJVhy9VL8NP/xf0UcObP9mc8+TDbxwZVhPnXlU
JWtS/E9e057+XWoO7ECY2HP65sDKuwE83jkT1xTikeh/7CsyEYtufMYTu+UCWsmGyXWonG1QM+XM
3ZmgSkua3KwnGE6nXsrXAbdfwR5WowCR+ld3+TYULHORFPZHu9CiLhri0sbUolS+44tYKhgbWyYM
0Oc/aOISFTcDmbEC5ucMk5ZF/uauBVig0xcigCqQwud2L0m23k/8sfiFdIjfgZw66oMojiK87Y8e
DfaxmnZZPuRHcSoAxx8pHUXctOO8THskIRpcxJkj02DyEVDL5Lu9FY8IaeB0w4kNvWYi1XgOQ1sz
ba0YO6mOqr/MQ2TTDtLrtNaOzRaPeNcMe589P/xYl1a62718RCkVYC8Zu3kOIYpl0hcadRurcS7F
hjGtgWFfIvUnK/xDmEXOCMrH5vu5lwj2CZXKZ9B063C/GoBEU4C6p/aveWe7530Nrx0AHkGo4nZz
utib/DY4i9jzU7QrCfnrl3tf3GGENUVrqUdFIQfF/bOR2O4YUg30zOWJHATiDOoved1ZFusz5jS0
IyfEeGxRJ/6py0pxcFqcyajATDlH7GsnplOmR+I61GYh9JLDdVzZKdnJR6LJ4vk3Cj69Es1zbX4t
AskyGmGuOuhVwf75K484cdROiz2orZuD3/U3lhW6M803/qyoqSYE3gz8Q+ADFiIq/ilLkQuJEdfw
b2aFbzVVMyv9S3IOB5r92jVOQe9wU2hazNr7abpCuEZWjIqBTmfuvP5LK6IE30qMzrYS+LNpI8BQ
aj6DNEJsr97z/iiqNJiNNTjtfh2uPl7Phjy05emTWOlHJCsD5wQP0VkBnXnO2WXH7nYAtE1YGHlX
2jK6rlLw6Mg8bJlIlEHHmc9l2TOGEcAaSVa69RyUlcO5tDl8TX12MyUkOL7ocwfrMqNaat8dfjta
hFQ7KocJ2ayL2scATo8kShIdllUWBZ4oS0IB1OhcSHnsvuJSt8i0KtdaPEc5/Vif9LMYZTwLU12y
MYIc3odweMiLCnVVikWCY2DEfqoh1wsRIalFgZb76bJQr8xSF056Gd/zOG34nGG+98VaYRacfQxt
2NQulft9YNZQH/Nns0LFhKhGqpPzAQtpHnEA79KLLDQ2jJeqN9R//nMBvzEGthNKzAqgN7cOx5Gk
/9uJKHjRsW3L24Pw/asPIqCqEMcdevaSPtB8g2HNZGu1x8NU+wrzW0O7PhO3qsP5iu4phP41j0ir
9AmduJQXR8m1MCnwo9e+LBgEtZnW1FqBiV0U5VquUWXrvnEkqXcws89iCuPuvlVPIHkJchofg+SF
ryI87lbrAFsEYS+JN5QKZujL1usNj3agFPkud+wJAIyyrTLIL5X5kxai/yVLiw6eKqEIbY1+qBNx
Gy+5BBjIRDEK33bFz0CpVhGLJs3h0cmRzJmIb5UNdFHjQq3EgiOnBOP/kf3MvU8Fxsn5AbMcOvXB
FaEUxjTINtz5Ua6n93U7VAKyzjgdjzLvaDrIlPJmw/9tX1/6bA2aUAIfhmzopderwO9OIlgb36Ab
0+1vdQ2kfHhDFDXeZ09Ea0bS+BZhZmmCxlr9acqPIdxFwCIuSFo5XXNlEl8PUddH39s7KrzbfH6c
JSlMJwsvUEw4eGiVtJWaDlCJ5J6/gPFPNCLcpPPOygfLQTPS9Pe6xHnJ9cGAWPtlWwh1iW0NmKD8
kWX3CjI74zCIcrmOq6f2FUp1IcXFbbxoE35A8L+rWovSGatpsl6YHeWnHvo=
`protect end_protected
