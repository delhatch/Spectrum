��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X.�84PT6s{W��Me��$�3��Y'o���c�lO����<y��CR�� �(V�d>>|��!��G���B����E]j:PhV2��	�x,�+�Ȅ0 w-y4���f���"I(�o���M��� �����p��; n
���ĩ�:�t�N]�Őw��)���t�k��xmU������N/��R���s�pH؆�p�,�wDo�f�k��Ĝ� :E���$�!D�F�Qj�%��܈v�k����}��8�~v;���:�GI�?�EAË�3k~I�M�s�� ��:���Pn������\l��1�k���DN�n�C��?�C��Nߘ�=\���������\��.ڪ�<zT.#��rj&)J2�����؛��V�
��7������ӯ�Lպ謋e=��t�m$(,��0�}���I﯄��͢�(;����߇��虵��}?��j;O�s�1s��a���V;)�|u3��}����u���a��e�ǎQ����OrNu�O�)^+\fHA!ϝkqm�RR�o�JPue�����]��e����/�y�C�d��5���~>6���l�0�R�禘�0��|�Ud�����������̥g�I/x������k�'�$��F�.넥�������8�?MYC�N7*�AWQѭY��å��Ҭ*ۑ�B6심��\�p� ��4߬E�Ţr�����`��@Fn���zcB.FZڷ�BP#��p��=��ۏ�!b�7#������cǒ���2Rk��D���i 1܊Z�-��.̽}���֝�Ryv-�-�k��k`�c��3M�ʨK���f?"_�8ZW�m�Ei}�-�s��ck?�A^��06W�MF
���U޵�5o��z��~D٭��}Gq������J�>rЊᇃ��v5�@�C-\���@��|l�}DZQ��k�v`ݖ�O�G\�Ki%�մM�J�"�`
�fI�d�9�OɸC�+CK�M�WG�H�N\��t������p�>n�0�����P�����aA���Y�=���"����K��s��0��x�qo��C��Z�c���aE�f�!�E�>m��>�A׵����4�ᓰ����C��Us�=��w�Z��I}�W#,L϶M�R�K�2L�}Lm��x�"Z�����R���c�|�S7� $Ƙ�C�_[��|����˽f/?���)S���sl�Ow���C_PmO'&S��Dqr�&�B4:%��1��Y�|�Y{��I����h��T��oo*4�̜�ș��p�$P��3o�8��ˌ�Y�����?&����J�]p �q���i����J���uX�刅��d�\�_
aB�?�p��� i�(��a���Q|�tV���d�G��dT4$Kz�!��s�T����9��6��&2rRUZa�7kdJ?3-�WJu��#� ����eaD���������C�xk��H%���\��[~�~�+��*��2ٖ'���6��:�nZ�u�ҽ�������e��4���u:ѩj��F,����1J��D1�m��c�/Ƶ$�)�jƜ�[󾏮إϣWYŸ����d����<���oRSڋd��ܑ�t�E��b�yv�2}�6=}���|(�k]maFRR
�{@��n���f�3=z��MS���=0ԯ$1�(��_V>eȤ���s���	59f_����<���j��Ы�$8{8L@��6�O�u�w~��]��-!c,�E,��gv���ˀ��:OY�J$��?�c��_��~`a�c�Sj|�y"_l�j��ք�(���u�#�A��oʂ���֗�M���!'tK㢁�ǈ6+�킣�$+�����TM�t���1=I��
��m�5i���p]����O�'e� ����x
-߂�^6�:z�ɺH��j��Y��S�f��)�N�$�>�]����&�A_*jp��!���I��Ɏ�K�2��z��f6�R��o��C�A%��n�o��Գ�4�"OܨX�F�P�g߇�}{��0M�8�����fr�����d�#��Rb��8x���*�R�P�{S�\{-�Wؘ�kp��.¬��$0k߈�mds�Hu]}���6�%��.ZNh<���&o� ޟ 'ʥ�N'+)��N����)ː���-�)1�Ӗ�)�X}�xs��y+�8�q$9�a:o$V�h�[�aY}�h���r0�Y��V�U��UL~
�[�k�Ci����߇�M�5�w��iy�Z"�Y�~��y�����16��K�aC-�9��$��3̱�w��BFu�K:	3�n��� �|�X5-и\�
{y$WP��w"�F*Cb�n�4e3����=�솦���Vv����-Jx��_N�۔4c�������>|�e��E ���9%�������S���Y60�c�*�d " ;�FO;1�[�v�R������> ��`ZC�z��m-��� ��t�7^�jm��벗���z�P�����沜N�.��Vc��>�>2�.=�d��wŶ�Ӻgf?i�"j����{�w����4D�i��_�~��>u9���뚿(աV	.�W]��> ���*���/s�6<S�T��{Uߥ�Ѡ������ Z ��cʹ d��h�̌l��A`�{�^o�wsc��L��musp�u׎�|Z��;"�b�b���f@F �G��T	^�s��>��MQV�t9��n�n���c(�tn�-ɤeW�"giz����)��������F�#{b�O��":�
�����%"n�|.�DY�_�PS�����L
ͻ�+:��վ�)�UPk%��Uܒ�ѥ�$�eO����5��!�X���g�ku��9��b,��oc�����S�%�']��v�I�k�"�P��K&�Ac�N���.rۿ�{R���:4ݾfv�Q{�٣��q�`�����ϴl� g�;�(��ΝRqC@2�^��4mQ�'����E-f��yQ�Zץv4��].�\�q#
��[!�g��ow@���Yq�� �G���}�e�_c"uv1���6�E"�����eh���03Lq�����S�NV)��	&�@['�[���ZR9�ד�m���x4��]�B<:^B�-�|�sA]QA�,�Y�����:�L�%�?M	uM��'�0W���_0�㶘i�W���p�a��?яK�qjb(�]Gz��j�4*�5�u�m��u�|,�=��Z"����a�5�|����|��%���2�_�"q?�_�x��a�)�-ro�L/�X�tp��D�n+��!�Y4����9��%�O[�c���&̓��8d�@_&ٛ�`c�4�lm��d,?f��My�_��������B�\�Zͽ�� ��6AP[`�9���,E�'�~��6���aNM�n���|@h�T��Gbڥ�$/��3%i�T��1��A����7�b�r����,�5+w�%�D���j���I�JVu���U����Ih�g|��<W�\qؒ��}���󩃒��9�až���:Jm2��9R�GJ_��WC�X<��;Pĥ5��@�С'Z��_�,�"���&�^�����Q�Y��Ǌ@�&�z���.��K�%��˒sd�����6�ŪYݟ=',�A4�-5�H凋F�e��EUN��y��+l���k�G�]�i1(��ʕ��n���K���\A���?���N
�GN���^����o�Cz�b��ϜP�h�-&B�6�m����s��Np�l��%���ޘ�^��H಑�mT��D�3������uP�E��Z���rR��wG.�l)�W�&�"�7D/s�֏�֩͌��T�ƴ� ԁ�<��ٹ�폿AQc�W�}��w�X���Su7�^4��J�rw�yU�2S��F��'����V���(}��ۮ���$7�և��������G�x���q�0�X����?��j˺��!��)�4.��ퟪ�?��'��1
Gp����r��.�����Tk���]0|]���i/왠=���Ȁ��r���ܫ��|�m��J&����o�U����*�z�R��W*ϭ��A�A��1���)���2��2�	�a4����g"�-'�Z���`@C����a�p��fu0�e��"E�.h�)��~T�ڋh�6���k��檱�I�"�{J��/%/����j��ک����ghk1�`��+��Y2%!��.R�
�x� ����l�G%~�Lg+L~o�H�2��{��n���a`X�Y��o{M�� 7���]H�=UD���
r�t�ӈ(3$+B���ɮ18ȊH�?��5�~��[�BqxFŚ��"���ϗ��(��`N^#9o?1K�rP	�s�ڬ��X ���M�f�`�vDD/LH�S������˾�=�+�)
�>��v �W{� |����'*} 4
RE�J��׷&��b���bӶ�V෿�};��
ʖ�9�7Y{�E��|VG�����[�����!�D����V=���͉K?1O��n�~��X��B�H��$��,��eA��К�Ii|������9j˰t�㯽��hs����D�SA��5g�B
q=��ȼ�T;ţQ9���#
$C�$������K�y��������ag���~0Z��IV�:5z<���8�L��ڔ���~�pqd?hg < .�p&�t|�y��z�mtQ���w�(�1f)Wj�� 5=bńfF�ۻ�F����x�c;7�S��	�sx�[��'jn��xw 9F|���K�YGK�jo�0�q;�B4�xfr疡��ѱD��<�X��,��E����~��O9Ku�#�i�	,B�܇��~��� ����Z ,w����W 
Cj�i"��ȇ։�ھ���;d�?�����NP�`t�f�c�Ε+�s�Q��K	.f��˒�E.�0R�5ZDcK�f����p:�r+���.�*\4�X��3lE���EGʿpM�8r/���������/����@������?�%��ĥi�� 
��7��uʻc���!����<݄���7fRU�;Q�~ڮ�Ј�dM:FhɠHw�w�gU�vWM��c"��c�舜he��g2h�1����[����J�+�&?!|m�n/��[%g�@ǡ��e����[��[�63�wIY����8������8�Z���;H����4kA���z����Tٮr�)"��!quy�6��_�xFB�ؿY�}.#Gog=Kj�"�*
�8ݣ-Јl&�M���(��3q�Q?w4q��Ӹ�D�7�-�[QVEZ��ȟT��{���1Z�=�Y���4:V	/Z҇�ʜ���چ�+��h�Q��ɧ�¬,T��������q��g^�L�]v���O	�lTn�1��s�Eg��K@�.�	�eJC�5IKg�1��5��7��p����|�g��u��盹���8˝���ӽY[ؾpFtw���-m�w��@��|H��D9�*����� �ؓ��MW={)2�n��~�n?Ud'q8��29(�)�|�TTa$ȓ��No��H8��"��ml�7m&-���;YLk�O���-b Y��;nx��}�9�~�dG�J�U�&JI�3�]�l��ΎzG�H�.����Mܪd�A�%9|�zp��N��a��x]M�Ye`��d��Ѷ,�W�V�74_,.M�%M|�Z.X�՞a���4��1V�h �??K�W0(n֑��#����u���l��0V��+>�)9-ARS� |����[;�����/�."eN����b�y����bi�_*
�1	�� �\��⧙�3fA������BH�9������B�O�=A��^�Z �ٌz�5X�����|E���QKvI����#�q���S]���wi�0zq?���!�����;�ٖW*�s�,�֣��6�5�j+����Dj�}tiQ��}�ۦ�����X%Y�4jp��C^��N�ˋ6�l+ӫ�r�Ɨ�"'3�F!#`^�� `b�C2AzkݍY��뭀k��'�kZ8����T� Wv���$r|��Դe�����&)N��}�����Y�7_{�(���[����B����)�c�'����B�jz+(��1$Ka3�!�{�sLH���A[a4>����q���ٹ��+jV �}��' ����v9\��J.����tͺ�mbRÀ )�Y�!�2�[�#�N�<���#}[�l��W����w�Y�}}��w��Z&���(vӭ��M"��J����t��ix<�
-
/�`�OJ�p� �*�pV�O��4��l���)��N)����v�А�+�}a��ܺI�ļ�!���.A����*�KgJ�CTf���J��k"����qѵ�Bc�*Mސ��-��Kx��?�3�6I�T��8�b[��,L��˯uq��k����b�ǡ��<w ��T�,2W.�ߊ���jav,��[�9((��`PQ!x�H�.s1�@��A��B2�zB�Me_G�p9#b�b)�'�,k;|�~�C�D$�?ɡN���LAV��tX��An�:��4L&�}6.�?j�T�9N�[y�_t0�k��dz#���1�F�kZ�D��N
b�ϭ�ըH�2��._|dz����`_/ؤ�)��4-� �KJ�z�>E�p��J��CT�K%�	Q�f�L5��3!Q0��Hf�s�_hB����0�(n-��[#'�7�-(
� ��Z���6��B�T�t+Nb�Y��mo����2�HV�+�X=�w(��~�㋁
8��sL�U�%�g�+�7�H��):�એH%�4�3֫�B?�1@!�7��<����*���uǬ1t��>T��y��r��2�젿��<UI���T��^:ɧq�7�gG�3bj���� �+�A���(+Qx�~C�����o�CaР�Y�j�'�Uh���f AV���{�:\AÛks~�P�S1Hss��\oo(��O�`����/���%a9=]�"�<� �v6I
�3�,�ԕ� ����:<�ka4^������fL7���L�4�)h���ܬ���cS@�,ϔ�3{��j ߿Y��(���05�a����Ë�bR�Ig���S�k�n�?0��͏TQ���<C��8��]avA���?�G�tw�G�w^M-Q�<𭔃
c*T���b&A���A�ka ���v�3�jb:SM0o�C_âe������k�-a�\#"<�kC8���e'���֗B��RM���O�XJi��t�+��Y0Gp����bP�8�A/?y 6$jƐ��å�A���]����%�/Ae�R5N��"W��4�דpm�p�o�G�'�!������:</� ��L��^9�D��RJ�ۑ.Pk���$�(v��V����kL��N;�W�{%��'G����iE �zC_%����\b�=Z7^�I_RQ�a�oW�ʿ)��`�w���Kbl�m%�K��S'1��������$����~�l{7mϮ�n�E���8��n3�H�pj���DW�P��ݕ�B��m �;���j�ÐN���-_����7جNz8L �ȡ��&�N6�Vd��c�tDCjsd��İ�S�\�Џ`��Ǉ��o��q��*�g��|���l��2��A��?��3܋2o�[���6EߕeƜ���*g�LnŬ�K:��>s#7L�m�a�����.l�(���T$��S%3�H;��z�N=|��nFb�j�6�^�r�䩅�: �����-�P���VQ���f��PU
 ø�|r��W�k{������6��������8/���Н���`��w�,�P�^�ڠc��79PtGj��r;)�B����!��ԧ���';��~V3�:}����Y��:zƂ��u�� 2��x����qq�TQ����Zo�o��?.ZD��1�����'־Ș"�L�aC��>�r�0���5��кo��cF� _c��*❎�cTQ"�N~Z>���B�_��"Z�Z�U��7��s=���.~�e)��~ma�y�0�6��:�gQ��
#H�o��ˠ*f׋��{(�x��(b����ԡ�qjK�G�����o�A�ف}�GvZX��y����ß)"��90b�<�v���+*�03�Fo�+�I�C�u����礦UX��k@aqt�׉�y�?(��4g����om�Aл�
7�xd@}�2���e^�KSk<Җ��W��A��8�@N���,窺�Rl[~+u��`�a	����{{�!f�#s8r뵯u��qS���`��ښ������}�Y�E�:6�P1'�{(����T�zn��w�:N�6����R\�&�������mse����&o˽��sA>/,i܍*�=������ס�d�)��"�A,/#@��`R|,"��/*�a�=�r����$8�����)\b�
K`�_q�G��'��:t���9J��S��gãW����^C�K�5�^��/@�-kų���V��(��m�Ob2���A�J�yu��;��$���(I�-�1(�k��M��nM�+Y�}�O �3����'�I���W��&d��
��N��&Bp{���g�FB���v��#��w�?��Lr��Fq�I~���U��L6}��}�b.ˆ�w����K�`$4?�6��\6.T��&����6ǯl��)j$Fu4��߾�dD�������-ZL�A4�+�n�4X 3�����m��]Qx�/�$�WdX����y��ūB�xj�������He��An���,�{����& �K�ǫJ��,�M���5�!y�;[�a�E|�j��y�QV8Ӫ�( �݀�D_���0���ʁ&
�^��:�p@i(D36*I��7-�(.�ؿ���^"g�E��C�C��Ej�g�^��>�[ ��Ó*��)�kY�A��'8��V���桲U� ��/W�������9[�t�B�*�dE���* Zs]+������Ĵ�p��ru�a��
S�v[ÿ&|����!'^nj�t�r���_�ʷR��y��\ɍO���7ފ�:�[��&_-W�K�Y7�[�ߴ���	�R��K���r����2`��W�\=�	tY@yO���w�ыI��6՛���/��W�A[�*ĭ� ��B<��$;"�*�_���eTe�R���)�_�-�a�=��Z��nȔ1���O<h+8��l<�����RΥ�er'����wŖ���遄�O�Lb�=|��ZT<��]O�E�4�1�Bz���$�LU}k�4��U.�)^�v�I:cF������Z���� �6D\~�-��ij�2Nӯ2����:��Q�jU�g����,���b&�L�=/n^�b�H���~L�QTab|.D����$<@�����;|���Q"�W���?U:|GA��-ϒ>(�hTh�j�!V��5�')�D#ң�o�"*�+�<��[���<�2ɪCx�o�@|�.����:�@��:�5�Z�ʓ3��=����R�RgFk�~?)?
΀(��'���w��)&9/;�C�1=��F���_���B��n���]\��u�N� ���=q�,:|<{zH�����M'N�=M��<��}E�C�zn+PJ��V�y���F�"w^)y���>܅�U���&��n��f��r�Q�C��*�R���!���A����pcһ�����4~?����7 ~�|��#$�F�"*
I�gut2�����>u�ۇl.-�U�a&�q9��@�BגpO�� f��>I�5��/�)^�i Cv���v�jw�D�l�c�����S҅ܮv3�u�<`�+�T��kIF�*��Ar��
�V~oǸբ���}�̣����YFKy��Hy�q�DﺘGԡ��[���Θ%	�ܯ8�ծ�߅EԳ��Ⱥ}�,Ae�Vׂ��;���T���Iۅ��4�s�|�X��M'jl�� v88�P���Q�?�(��>NbS0,��X�A�ŠVf[����F��NE罣s�<1�7���ׁ�+���Y��)��]��Q���uO���t��`�.꩝>z��0 G�i�X�b���ɳ�z�[�a�h��������H��@���N��>��BcA�^�b	m��;
{�e�lA$�7Y�^���.��q�U���J��T�V�vٴ�|o�j��b����u�t%lk��*��i��� 16["a��Q��K5������)9��F&��hH��	{�zK�Cĺ�x�!�W(�ҠT+��nz�k��슍�]5����|��f�u���XR3���q{�0+��JS��pV=�XMU��B�H�d�ś��	�?�Pls��@�����}�߇����ϓ|�S����=��-0�e�Q|��A�1c����	P�Un�
���'��F��av5�������0/Lk�$�nZ<����0p��!��d5�{A���4��i�a]��3�8L%Ե���+�Se@��ߣ>�����'��`���G�.�,�ͿLᵳC~����N���x�B���7h��1��Za����ޖ�1@ث�r� �9��[��H��0H�I��{��ߛP?ؼC9�E9�"C<c������Yω��uQ٤��.�6�r�A�g�v�l ��s���s�!׫զ��#`sꖃ!E7��N�D��0+)�=u702�?�ԅG9#����/�^��D�>�f"��w���^�l��Å�㵨h?�4h�<���
�F��:�C(����B����w�ʘ��Z��O�Fk�\t��+��\�ʶ>�wC_ j���d���`D'�q����l{ʄ�S��ce�(�c�y��}�lE1|�&�Q4od~�<396���B�5c�b,-�d�(�?�J�d�V�ŷ�x)�pއ�������$67	wI^�h\���.g���.u� �Cr_�Y��u(#�d�*d�2q^�k��-��\z��ܣ�~���ŧvͶ-4?r��MI	vt\�G?jm�����#���e���}IT��C1e�"��Os��Z�7(	J�݋�Vj;U��hŊ�=�$��&12�2��no�������o�{+[�Q9^x�n��\� ���iQ�hG#)��ѼK4��9�>H�P���j!���-V79�$���:Y���f��Q�\��k���XΏ�m��X��g�LDӱB�d�Z��}��N}�s��V��mQ��]�ҭ���K������u;�~c@c����\;Y�q!�3I�R!!���܅N��%+sU~X!����Ac!�*6�y���B���IC�7�}�>�>m ����}��Q3�\�0�#��n}�F��v�����w�*�>�1���l�k�����PCj�g}�0�w�{�F�'I�fMW8ýL7*��R��_I��� *i	Cizr���򅨪��{�������b*	>���r�B�Dc�ٕ�rh�$�t0�rK��e������o_3��z��p��eG�6�����4޿��"I�n���Ī�E�
1�t�"uGOB9�숱p,�P�/�c�]?���K�m�u���&����V4�*'}J����j�w��
����� U'JZ�9w����WDE O�[e����U�HL�ީH��@x��]z͖��{װ�N�jP��yf���ۙ��]3D��%*�}pY~�7a���k��l.�Sb	s��g�Kj�!��j]
���G�CkY�¦\�%��!p��0d���.5Jz#��,�bG����o�q���ێ嶧c[MɭU�O�r�
�	a�dX����4h�0��nG�����{֓�,G���5	�O���JQْ��]�|�qr�C@�yX/�gY��$��C�޸Y:<�9��m��NF�P$�vuQ�(,��6ī���h�>�3s�$y��U�z�OH-��.��4�7M���V���h0������/�����,�0O �͔�o�궰��b��is1ʩ<�oL�>X�<�n(��zO�$��8K��ɠ��/��� �{Ό�<%�h����a�#���@v��U�p�Nl�aOxJ"�B�~�u�`��+8�
������|��;�VyM���L����Q�_ص�i#7W��Ŧw�i3��<'TQ�(#���I���d��v���eeIѨ�ZB~F�"�r����mCH1�0����L�;cbQwz�"sS��C1�D��R���'8��|d�+I��7����\M4�<o�Ge��Cr.���u�{�:@m������ɬ����<��Cpi�Y�8<�@���m=NU�χ��}; �@H��B���j��ؚϣ�]�Ǹ�v�/�K�1����<��م'g�����F6��QC����%|��\-��޵�ŊV��v�-j�D��$�	�
���-1�ȱ���I��v��=J�ϱ�c}��Qp���&����\m���ڧ�`�h�x�NAa�u���!���|��F2�����ٜҽ�.��e�#f�V^壤��`�Y�g�c;�� Y>?V�L�m���N �A�j��[��Wz�n�7��K��ҾG�dw�vJ�2���]�����AN���C(�.s�љ��a\�����RϹ�B��¹$�H)qSB�X��gv�[�JR�{ĥ�7�׸�i���l�^Лg��S��v#��qL��� ���׫�](�G֨ؑ� }�S���7)*ԪX���2mxw���y\��;Gri�^rIr��QC)�[ɦ��k�I �f����ԍp�5xgS�:o���BjY�y����75��R@XJ�'��=��Îrk������_yk����&���c�H���Z|O���l��:5�42��|���I@��-]�˔\_:�U�_ƨ�0�:t�.D�0�w��NREmnfsl��b��"A/�Ѓw�4��V�=���ի�'��hwJm̵K��:��}��ؒGrHYJ/6Bo\[*������w0Q���z9�#?Ew� ��UV/�1GãN�b�P�v�N>|��t�bu4�32�ʶ�J��o��>ɝF�jA�I��r7d_ؼȅ�����S]�=�<����9=�}ٽ�l�A#H��cz��5����f������֠�C���4�F����v�X�����h�=q,�]�*5Z�A�$G�-�l �]Y�b>��jQ����|[YJz�lmKT0�蛯@�^\��y�̷��ҩ�> ���IɃ�y�U�M�]��>(��Wjf)S;��2�q؝��FJ-ӂ-��7O]X^;�j�Ӓ�HShF��*�VlH\����Fy�A�4���k�FN�I9�{ҁ�k[[� me#a�l4#����~|��Iy�~����%��(���q��z�	�>�����K�ѻ�u�n��2����|T<׮Y�; Y����Z�:f�#���^|6/1�@��M��X�Ǟ��A��(}y�+\�5�p)��k�]l�u�y�(�ci���.�����4ef/H0/HSܧRT�8yY
ۚk�b������o+�}P��d-���Bu戣xI�\$����dR��X�}P���5�@U���I��A��)��
�]�J��`2��R;źN�l�g^��AM M�dE��~P��S��� ӷnF�Pڢ�H�a��":{�;��5۩�aW��=���&dc�h�-tciNA�F������>��W���:tÝ�n.��7�ihދųJ]j�JCwd�ۯ���,�_
H���C3�c
�"��W����=B��������@�֔� *�+�k�r��0����(��Z'��n�}ZT�:Z�|�:�r[�������"0�15�h�}�v�i�*K���8�M������7�b�bU�li��������)��c`_�����@@���3�1d�-�I���^�dW���tG���!<�8�D;s��ϲ[�">����CB�A�1k,t�7������?�G�
��:�B�~�l�E3�L'�0�S{ї��$v3F�.��"�Je���"�R�g�����
�nݰ�~�(Ʉ�d:Kt���-ҍq7�Y�2���نS��L��ܸh9~�+J�W��:ttidٟ�^?���8����Cr�סN�'zb���J�K�BU�=Z4�Ɨ�j�?����F)�*����Yi�?�DF�b��y��mj���=}c�M
#��-��"�"$ZS_fui�7I��hP	�xє�Y<��ב-���ȸ��j��Xp�H"��I^��� �'������r�o��0�*c��B��K�J3�x5Z�t}�)�;�p��ʹ@] Pf�7�Jqn .K钌�����M��/qЃ٫����9��U׭�@SR��
K�������.�P�>����	��l[ei����2��x�y���t���־���?�=�lZl+�[�<G�����'H��I���R�y��2sp尣�o�IL�we1Y練T��OP�Ţ�$�F��H�mJu����#�O�o�b���2v������ɬ�u���=�&3'��!��k�MEЉ]��w�i���y%.@*̴�ߝ���3����#t�c�]�Ͻ��uz�n��a�*3)�s<�hm"%60�0IP��>4CJ�EQ�H�K����j��v�V� ��c`�[
a^(�Uɝ�A\��-���4v�ݎ��O�"v�6 l���^DrD5�&y�H������r�~�p/ȥ��cZ���f�h䭍�)i�����g%�����,�l�e��-�[(�\�3���bZ�S!��U��ױ�D�s������������~;�D��djZ�T�.���;����mr-IM�E��m�\ju�դ"�s����Z0�ɇ*���"
�ͩ9x�*9\�����O~�z����_�@�$?z�]����h�.�b��w��;e����Y������>����l��ϖ��tЈr}P�&1v�{�W�!T�����̨/�Y;�ұ�!j��>�غ��Z!S���s�eI�31����鷈-'�ds?C�D�|s9�h�F�Z5kĶw�͎ګ3"Д���I��#sV]G��Qu]/�(Fj�r?i��h�,�r��� �����]r ��m��1�Ӎ_>��<�	�ٿ�ù
94=uC�7>{�@㼰�/<2���|��,{�U����'O���3���
�B����ME��0���u���V���ز�eL<��2�>ֳ��xWq��
�K�K��<L/ЧB�dҨ���ɱ�U��ئ��3��T|D@K��E�R��tF��`F�ֳ�>�-j"3?��O�<�	S']�J�u-?��M�<>��{t�/����䣍�"��������Bgܪ�~x .pe��k����S]���6��ʔ�	èQ'��5��%�9��c�)BB$:�&Q�����>k�`����fj�"�4n���ԶĖt�}TL����_;r� |��P�q?�ai��BQ�C��ȇ��]�V@�3r��g��G�Nm)��>�bI�B��7r�_ W��60* ~- $�uд6h�<��1\=K�Vl>�1��Ch�(�D��LG����`Kh�;л����$2�"�(S)4틬��1�vuj2���!b��[`���n��p��S|���B3��#�y�1�t��95,YR�8_�x���'Yn��Z�?�n5z�`P�����.�h��W����+��;@��6)Tg�#�(��x��TG�f7Բ_(i2�M�]u������Z���i��`a�A��6d�ӻ{�YC4=�p@�єn̗ʰ^G���\��u#8c�]Bf�`&v/h���5����s�z�����o���k[�leF$1��\�m�6��O`p�]�B��F��j�����[��ӗ[�\�PV�R^��>���e?��r/J��If��xT��é�CW�e��E�\>R�ꀽj]u��R�Ì�8_'<u���k<��^�u��f��a�NQKcy��W�%�$�1�j�B�#e��1��/�9R�eqLt\�3��I�l���*A2��n�^��"��f���R�M����c��䤳�7WhSnUع�L8/˩��>Q���]�e����!����h��m��~����~�=�*Nrqf�L�K�����漙,u�9��<���;��̈qH�ґ�3�z�Y��Y�
gu�d=sLF�t��h�/�)람'D\�Rɿ�Yɉ��}K�@�v(�eW�ݳ���7������x���
�i!Y�l��� M��|`�6%��u��ۗI������+�y ���c#�ːpc����oA�Y���R6�P���+En�Ӱ���Q��[)'�P������%s�]Z?������}�[T!IS��tY�ַ�6�Ͷ��=u9�$Õ��z_�p͊E�ilj��ZѠ�IzDF�D�3��y�x�d�������u���X\)kE��r��@��=D�����!LF��Xu5�v���/�K������:0����xWQ�\��L�E�c_FW3���g��| ]6eh�
�y9�QpW2�2GBRKaG���Z�,�G��C�E�~���<���U�%�)���i�3-ҔM_�|u�˓i瘙*'�T*�ǵ�w��z'&a�/:�\�2߉�EFo{�����*��0lG���ɣi{x��~�8�@��[*��MY��Gh .�@|Co��i�GE���k�
L�і����a34���Ȍ��.&�̒J�Y�z����AWE�L�$b9@kxn	�rjX
ˎA��鈜��Ѓa�S��a��'��U)"��dՀ�a�]jF(Dݤm�Q<�:�e� �~�f�W[\��Ayıe�T[)K�SQ�{�T�� >�d�2�_�r��1l �Z�S��d�[�7���˂P��Z3��g�(��<Δ��=�c��A�.����J-�Kd�*YJ��ec�����6r]>b1Q�/���b��2$֖� 
�����+?�D��oH�k��낌�'� �Q|߭�;w����� W��!i�
\ғ�î���_)u�o^U�dg�p#�^r�ruw�2���Ѓ#�w���+���&��X;BV'���<!d�b+jAj�� Yd��9�r=���.T�eG?2��lh�[Ĺ�/r@�=h�|�գS}:)��}噌(���l��Tv�A9��}���ʠ�&�om�QsJj�@�"tZ�6�g�
l��� �u~9�6LD���:���#��m4��;���0�#���dK�L�|��TJ�w��f	��Keq�ϳ�d#�/o�4��y$���o�㤩ig�+�2� �MH��:��_�a�@��&��)�18C�ؽ(T\%���h�7��9��ٻ�U��|=5��_�d��d�khd�h2&��[,��^���9��4aB|(�/k�z���p2��\��$1��ǎn/*\� ���_P�����b�ў��4��S�ֵ��q�X�l�T4hJ�^���Xh<�M��Am�L���:���S���:���Ӌ�g�x	�0b����������&�Z�P�.�,.a3e��p@���2��Q?�&<�����*�j؜��dje�w��i�vT�x�,�#���5xe3�3Ri����ҷ��&S�&���^��� J4���"�{����.v|��Z>��E+����"_��׭,��*n�'�eznŒD�T�|e2�u#W3wd�9�e��L�&���a���U=L�y4)���~�<$��l�Q��k�,�@c�`����~��xOk\`�����id	kȴ��L�X�s��O�ݻSΨzJ_�;�9^����|�mڱM�|�p`Zz&˼�~q�\��8-z��'���L1��s�1j��bUvC� Y��1H��|�U�+uE�|���B�����B�x����M�Ҥ�*˘QԆ�_�����Pվ��Ro�]D�IT}.t_B��z\���?�����{��(4b�e���f����%�'�9s����ƍ��(T��[��X�N��-MyP@��1f4̒�py䁻�`i� .Թ]������@�W+-��@M�\L���M<��ڲ�A"um�'W#���9�T�K��<��ǜ�S.eD��l�	1I��5m�̤�������6���$�e���j̾����T{�goͲ�l���B�ub�`we��n{;��k+}���;��	�^�V�e�q�N̸Ώ��0�XU���k h^.Z�#�Yҩ�o�cr��s��ؘ�����5��L��f0jX<~G������Y�uj~�{�f �C�R������~�(����׺����D��-89lp�m��`���}��>1ti��6h�6���oX����_�)�̡�_�������P9- �h�O�4j�>Hj`�jT,a�ЫTf���Ń���"�Ϭn�]Y�\?{�`�x��i��gۙ�to���lHA�.n��F��̭��v���-���E�{���Z>�yU�ޣb�*�TL���v�7'lp�}4�睸��&Ac� �js.���&��g�+�R�g8���݃ii�hl�{�߉oe�0�Q������F2�������b8���B2��'�����%#�W���*�AYh�r5=W���:D:��j�x {2��h����Z�.U<~�u�1�G�ۃ��DԸ9v�����z�x-,F�vu��*(��A&���.��ݓ
�;�݆�7�����t����n
��Fȃ&.��Nh��m��A�������q�t����с��ף����￝;] sk���;���/���+8D�#V��&T�v9QRRUwǝ.Gn(�g��"�u��B&��������l�Ć�x5���'�<o�Sؕ��qQ�WE?�5!�e��h�'�#1a���6��w�a�u��~�c��ɲ5%i���#4~������Re�=�5���#6��Pd5�/#h4�ǯ�T�x�.?�\?���zq��ua��	����ypގ|�}��[�4�-}
�.���x�N���!I�#�k����v��8�ڵ�4�rD��#h���aPM�qhv�MJ�88Ȁ̸��U��ih���C�h�=^$�1�,e���t��b'�>=Z%		��0Ʒ:S*D��𠟄)<N�-ܯ����
ܿ��������>Y�c����Ŧuw�+�t��,��j����}(þ��p���1�;5�3y��zO��5�΃�y�Ra��s�E�|���+>���1sl�4��s��B!�O�wT�lph88�~�
'�ڨL���~9����k�,Y?#��ooO��� ��2"{�A~ҵ��������u���~ЩJu�仟���0ex��
�o��k
a�ao|f!�����:y�)ָ�y�W��zc����(g�2i��p7⻵�.��-����1��uY|�Z��|Q[��9�@L���A06��H	:��e�9caI����
FQ�Fc���e�q��<�7��!�f&D�ɣ�X�+���~���3��4`YA���P��6�QX='܏��Dr�B/3�t��v�����4.]_�d��i�{^*�A���G���-w
KZ	�'��̕��T5q��q�OW`{E��tQG9������ �=��X�+i��
���d��}����p,��������n��I����X�la����_�-�Ad	�+���G1�� u�{��#�O$����D
����p�a���س�^�1q�V�#�mZTѺ���,�g��M�efZ._:/��_Ϝ�y�ރW抍T�����N�}�q�b�O$&��6�]��i�iZ�}F�I�I�uf�������#,���ы�]t߯q-C��D�ؠm����.����@�'���H�7��i]�P��@Q���54qh��g�)�-YBmq3�X۟�({�2���+� 겗 �~,��h��S��;��؎(DzX)�2��u1w�|��ç�f�ʍ.(�d$>�j����7��mmi���7�_���5�2~(
����?_�h�)�*,�K/��ή���\B�!p)'�p���s�3ҩ�r^���)En��M�o]��3w�^�A�z�e��өc��� 62'9�s�A�tR�Nq��L6d3�f�q�R7N�>����K���W�gPp~K�?E���&
��ɔ~v��Zf 689�G��4 ���~!e6��z,��n ֿ� ,0{��\��L,��dOT�&�^O��^�C�4n��\���/�Op2��`e��^�=�b��Qe��ԵK�@�Y]h���������X���tō��ux'BD�ǤRS%���[��r�3�x�Ǫr]��*�=�PΧS��Y�����4~�� ¿2@�_��N����/�G�0o�2��״E�IC�S�p{N�$�)�����I�;�$���U8ni�^4���T�D<�bL��pl_%��g�0���3�s�=�s��`������t���v�$q�>mq{�F$����wF�[�����qc�Ew�2j���Kl��cO_���#^I%�P��'P��H���a� Yo�Ȭ�(�噀Z�8��A:"lnB���c!8+Hz@B���m?c�Q�q	���J�����v�����d0�֊�� �λ��>��9o��:3�ϻ�Q��R���f�c�'��m�	}K�XGD#%u���Yw�e{A�i��g��)q��cQÛ��D�_N��*�����WS�*���O��Yr)E[S��ݕp��I;��u��k�)\Gڎ6�3⅒H���)E�ڧ��9��M��28��w�����w��7��:,�z�Q�I�p<:4�Gg3vJ�RI�&���aa��VB��d�Fxwt�2�׫8Ԩ`vcb�|3HAP�xa?��� �������B�h�y�e$��VT<Ԋ��qGnL����*������a}�B�`�H��$Â0���~�T���N+Ӱ�(�J�:yb����rpMҖ�%��*&Ϋ�% X�pVX��y\ƺ���".��e��@0ё(<� ��o����rVDevk��Ê�|��4��7�+����	$Z�X������`*\ \UP���>A�{�q�{�C�A9{k�ã�x&����O���j<|��G�����怪2d's���Og�U�Iw�ѐ"�{�qH��}��P�9h�mi~
g�X��Ҭ$T>�8H8�r�������b�n���������v�Z�W��-Ca���I������S��N�7��m`��I����a&�4�4�X���~�7?=CD���A�����,��m��s��l�j��i�.�����.��t�qm����$O�(&�dO��A�I����<�c[�
�������M�ࡍ+NxĠ.�/Sd�H��:�rb\�X3�V�2���`�C��}�Eo���y#��5�:�-��h�t�:�PT'H*�6X<L��^$�7�>���