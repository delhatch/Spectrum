��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X���r��Иwd��G�<�
�h0Jj���%��ݜ�.�D�=�7�_D��~�~N$�o�0{��2�2�Y�����NSØ�?����k����KNlu��vZW[���$�Ȩ�V)�5i�ӽ�DNkev4����j�Z;�8�{E?tȇ���f��	�8�w���gX°F����rҠP�@���t�ܠ��Ιg�1�וҦC�}�H⍌qv��K��	d��u��Y`2��?��ORn�� O�E=0��H�h�KfH���␑��X��R���wl!)k6�ܢ*9�a����:w��䆙�S4+w�������/v0<0�c��p���Cmc1�;����VV6Y?X�cd�����x཭=��=���ͣ�Ua�L?���˭�r>o�w��4k!�eTe�J\�����T�R� �Y�}Zn5���q
Z=��r0�b��D;�r���)�?0� K�p�s?>�|؆M"P�3 �R�0~�v��2?~��-vɨ��������i�g���u��� K	5�Qܱ��M'���B����K��΃�`ٵ�0* Z��f��Yd�7����3�¬���
F!�k0u��<);�R�J����=� �SQT��<�0���T0|Z��ư�XI/Z�M�e����K�O��,GZ˗L� ]'#���'7�{$������0���"��Q����l�ceAh,8��?���9��*b)��ˋpӰ�iA��T�,H_�]d��R�i3�:��6��d�
���JX$]�<�Ģ��c\�W���$�ߕ��x�Nz�b�A,Em����)�h�:G���P���)���X�����੊y���T̹Q�x���*G/���Ȅ7M}FH���頁 �hw�}W�2ܥh����#�o��ʱ�QG(�O��U�Es��W�頻%�)�G���O30�S\�����3W:���."-��53�Vk)���!�+��DxX��D��1ⅲ�d1�F!�R�������d�]fIT,��!FX����u�!�[����l6ڐ��\g�LMW�R�s>uy�rk����ğ<w��VJ!����{�s}L�q%EAz#kIdOM�:��:2ZS�h�o[pz �9�ӂ ���:���EV>��(m��FJ��ɞ�Uoy_� _F�1ь�<��\�䮀b��99q]�����B����Sj��\_X����HY{�"�3lT:lǭ Q�w����;���t�`ȝ�R�)�Oz|��wZ8��K��;�ԇ2��������g$G#6u0B�@=(0��k�G�w��|U�G���������.Мe�0,�a��5Մ^ɣۖ�*vX�
K���/\&x�)a��}�MOs_lYj�3�M�k�ū�F�P�f�Za/��l3�����`�h@�%.�v��P������n�ߩKM�N�Mf&y�o�B�81-�c$C��^��9$J����?�F�'�/؎��� ���'#��~�N�~K"�@�8�?W_͞����I۩5��˪��cT�x�QF��$x�]���mltڜ�� ���#�VP;X� ��?&��H��5�e��^A����FRv�D��:睊��r@Ƀ�V��KJ�C���I�$[�ġ��,��3�Vf|M�׏q��E�E�_��'5S/���ʍ��n)Y�(,������XxI��)�.V7��
��P�6n���n�S�Ň}l�X�<���*�ᙣ�~p!5PL.(�f���*�-�$L팷7�0�i1�:�[��+�N.\�[-W���Zݰ}�v旸.�%^�}2a8֐�n���pU��V��B��CB�bv�k[nt�$@l��(��fWN�̳��>?!K��)}|�Sg�ךX��2����l��[��wr���������b�����B4A����Q�u�ܦiM���-n��胹��l��9�L�"��y�+`S��=�����V@������BI�����-)��}[�'�༿�Xa�p��n9#%�R贑M�s	S��k��1%Ѷ�8�:�Nm�R���(�T�H��#��N�H,�T�Fkͪ{]oc�r9����yw�Մ{��������? �P��p��tW�W��-��/+u1��KP�ttm�H�zUv��]z$����*�?�+���v<nB]%o�b���ڂ���J���Q��Ѓ/�Z��F�T�#t�oL�}5Y�8�I�[j؃�h�-���4�0{ښ�������|�{�τu9�E&�xh
�G}�\�D�c4zog�Ju(ô2��>�ttZ
���'��&C �,��&f��ٴ��%�!�)��<��M�d���%�ѯa罬��V�"�+���[b��,�!(���34��u���}r%�Sâ[�<O_.sOt�k�h��DZ��їiL��6�i)���EC�=��7T���z.g�$������7�K�m��K���Zk�YU��m�~�X���ICOGo$b$�J]a�7�ny��~����/����JT�L�&^�>B��.)/x���׳���:ܒ�� W��%��O�f�ek�G%36R慺~���:%՝&az|#
�ʆ� ����[�+s��l�H���%bf�^�A��ɂ2W�Zm��:���2YI�}�U�W �t�,?M�W|@M�g
y�p��b�����U����4��$):��~?�\�c��iv�<dDh��-bbM� �T�k��C�a��m�.��P��q��!R쒝i�^�l��ɜ�R.g�&�&���r�{I<1�i�gJv�K1��s"hZ�
����P_��:��
'��u(iw�Ity;=����8��rȐ����aHfۦʉ;��e��'}hrj!��
��� �u��:�Y�hﭖ��Y��4��%�ʈ� �h �a��G���3||����A����3�͛F�؂2�(rz��r͌��؟��$�>[::2kr��HcB�b�0��z��3�(;AR`��y9*�?�Q�&�"��)�ۅ*h<#�ba��K��j�B��}q�jaT�V�'r���u���I8SaB�m�� c�ik�_(�#��[�� �GFd�����UL�e� �[�%_GO����R���N��a���Q���j$���#�wdh��'ߑ�<���{b���Ӂg��^��1SV�;����	ۆH����=ˍ�9]No>��!��[N��OY͞n��y�n��6.�g���'�\���u2��&Zw��
����_�nLA� ���0ӕdL&����v��,F��F?F_Ԯ&��j�o�
O�b�F";��?{u@RU�E�p���P����Wl>e�8�H�V�����kД�B;�@��"��!���3�X����xp,%l��\�V3w:�L���_Kv~��r�.(ЪL$�R�1g�;f�:�5>+6#�:��R���I�����W�N<��� eq��d��V0���?@�L��ٹ$9W̺>���'���ӰH��<���et_<�^�PQ+���i2R��px6wG�_��7~����aR��i-	V���5�X,5����Q=�ªW;CL�%"�1�C	�4u����e �Īyi{17��v��������Z�:DQ�g�Ŧ��r��*뚷�ޤ[G`mZ"7RJ�Q`w}�}�@�<���S�@�q��׻ɬK����fq��h�3�ܸ�J>�dZ%�#��I�_@w�) +��k"n�5��l������s*�7���D�y�W��:`�m�C�����.�^�ɀh�Q���<��6��e�eE/�B��1��&��;��,2�?g6O}Z��E��)�����^/�ZA Y���YB�$!�}�ʲi�;ު�|ӟϷ��};��}.�~�nd+D�H��m��s��{��U�PK���n��W�,q؆�Êu���W����d��Q=�}mb2/�z'y��J�0�3�<pʲ^�I��2�7��9�S��
���uc����_8[/��'��&���d#ǆڦ���$@YP����<�d����Y��R���w�g>S��o���I�bq��*C��TPFʐ�'�3�)���z�XY�~L,�q(&[{i���k��:�*��+\�c�^�t�I3X৘*�CE��:�q�I���r��G��-���!��C����U�����3� ��Tuk3
u���|ƿ�O�������?���ԵZ���>� #iu>���2*�^�j���	���7,N(l���y!˱ʦ���N�d�C��Z -r��/��T�lҒjx[J1)�scsvQ ����2��1�c2>w���)' ���Ra�w�Xz��=\���J��Kg�?��;�S������ʛ���Ҽ�B/6�:_��=Z�P��4G��
���x�9�n1���8�q�Z�$iQz�㑙HNU|Q�c8�&YK�k;Z�%X7Sm��a:���`����u�', �!�*�<���e�V���0(Կ���N\������o&.<���t��?>�"$�͌�GP�e��w�FG�������|���;Z�ݤ@�b��V�׀g��H�&��f�J+����������׊S^;�=t�U&z�����q�/v`��#C����_��_5�80�?O�'�1��޽%N��4���Y����^瑸���\�6�7[��|C��VL5��.�'�����R����lԺ���l;^uf��I01�P�͑��#����lW�q�x`�Y��L��4(�N<��6DP��Rw�Dͽ�PӦ�n��a�!�O�E ����޹n��vck���a�Q�C��o�%o�|z�
�F��`p���6D��:��d��ݥk!}�@2���_�	�pb�@�Öw �y&��Z0�� %�}���X��W�X;<S{�#K�����^.m�.���0�.���6<M��{R2�0�0<�	 �߿��W�e]n�f��(��b7�����Lc���/嶲����:���c5��вEN7����au�yZD�b'��/��М#ڽwB���U�Xw���ٱ���Y���7��]ͧ�{(��D�U�j���d+��H|�&J�����c�=j;��(�N��(�<�RB�C;&f���}�@�Հ�����̗�d���.Np��)�����oP����`� ��2$�����VQ+J���)W0^������!V���3�*,�C�B�(�?ū/&4O��g�>�3�},{��G�J	��ѩ��RT�-��b�]�A�*5��o����I�a�YTX}5�HQ]�i���͂����rX\N�|��/�u!��r����٭D,�� $ڽ��N]!I�/��\��X{&x�ܚ�M��%�ۜ�;,�E�]K���R���t�t��Dj��
����N�g�!2����I���<�	�3f;Qg�w����/	�8�w=^Հ-���-��^��0�Ů�)�4»������kA�Cç9x.�1_�*"�t���sFh��
Cͨ�LN�!R���E���c{B�����XFpG��>c�k��_z7ĎF� ��|O)�9ڼ�b֟�0��%��0zu�˦>PF�<.�dR�ئ�ޜTl���q�C�\zL��B�=�]d����yN_�o��}�VC�������ټ�O#��_nkx�κ�*��Hnq�Lg�赩��:q��+�ښ�h�mk@b�9"<�i&ق�v��nkf�܃
\T.Њ@���퀔���_���.�2q��:�j#����pE�`���;=�~�#b��@6)mTRt��n`3��Js���I%���7b���=�?C��b֕��[%�P�5�XW����'������`7��N}���>t�?���b�����C���L�h-$\x"�/���g~Zƛ�sd���1;�A��b���vj�ˉ�����ˣ�X_~�>�7b��M�Њ9��mY�@,�]\�� nd"S�$��u{�����v�q��@��4a!�>�3�A�]<Ŏ�"��j�X�e��!&�ѷIj�qs��T����<��gW�˿���y`�]���u�jS$�k����Q�\fU8�=0'�1����!/����:�np);��B"09`F��Qy�|��3��91�2.z��y����43D�?޽�;�R�[g<1<�8 S�%�|6�F���)�T=�R)|�W���� ?��F��d*�1�Z��`&��C�cr}��f7�d�C�;V�>�Cr��7��bjus�<�y�)xY��+���M�)�!����Y�O��A�-
b�L�PK�xP��e�$����]�Q^h?&m��T�̬�b��\�W������^C4�ʧ�|\V���#����cÇ�7�-���y �2�٫Ώ�Mg8iOhl9���r{@�Aka���N�KXsv���ZOК�z%�S>�R���o���:���R��*xN���Gu+=G�>zX�P7xCﶺ$��������^�F53۾���]*2wH����.+0����������xLdҭ���oK������M���x`Ţ�_��̃<G�ݹ^{�IT��*-8��/Mz�@G��
�� Q�<��B��#���[�wX�Ќ)-�0	�(�Q��@
�s/j������֥$�����Ӳ;���+z[�_��@��VV6��Mb�� ����bN�il{�7�_�N��Hd<8��W����^���q�|A��QL d�kg���xO<��#7��)�Xc��F3�^�M���u��W�l����A�W�<�&��k/� %��Z6���k+T�Jإ��H�zY���;j∣GmAH-�{\'NS��8Ķ�V&���4�
��[��fU3Q��&��wī��RvZ�w��Tp{L_��|p;dK2w��7F���_��v��=ړp���<�p��ex�HRj�!h��ͣ��|����=j�.ܸ����s�����!��_����<{7�S� �J�y�b�o�6��A$S%���߂uiɦ1�`��ˊ�RȄ��[����*���%ya������M���K� ���%g�mۀ�4�T�&��s6����d��/aη�|�����ײ�uTe|��I;n�?h>�`x*��2'��V����#&T�;��w��M�V�
�=.��)UL@3"t��N��{�Q�{���E�|�R���.�ʔ��PO�É��R��P����-\S񈞇�t.
�/r� �8���q��i�E��8�g8)i�M�RP�&�:���M���=cp�H[+(�F�4Qvt9�E;�i��?P�f[�/���p)K�;��Z�?rpR:K���򌻠~	�H� ���[�q���S�ݳB��9���2�%R������B�o{*V��Qd�9��N�:b&"2�;݆a�]k����8�,|=�; Cӣ��bB9���0/�w��L*�ۢ��{�e��c�&:�!u:�l�l�̀:8���9I ���zAk:�^� ���.��8G]��O���<���VH��=Z��A5�Ť��"`����&�/�);��0��NG b93��#��s�c@z$�}�TL�/���!����[cO��s��=���,-�>�m8�����zD�`$9�#���:��Y��6����@'\��h��'����*p�m�7��>Ƥ�Z����
��Mk4Pv�>�2w߲_���;4��r��L���o=!�W���{qe�@t$�Qf���{�hsd���W5d�f�s8X.!���*�T�,SfA���d#H�����6��^l4OwZ����t��h\doB��kM���v�m(���:���'�a�␄~ �$��߹�o�U�kY��ҷ����=[0�1�!��!�P̓���2��M�d��5:�Qy���@}���o���05��|�4��=�y C��Z ��q�O�6O8Ó��ňt�8|��	�}t�2�(5Q��y)QO�+��圜����ajނ/ �<�Y�*L(���=S8�lM��q$��L�Cj��ho:�`������.?B�����a�VY�5��b��}91V�]�V�Jx�Nja	3�y�D��SYBM��Ͳ�tq*����f�+�g���4&���!/yUHL�h���G����gI� �k$�Q��F�j��zE-�+�M��p/V�L�8$�V�4*@o�0rP}]�r�.b�DNg���~A�wŉjw��+ â_hᭇy*ŏrS��m��v��<�Q>sQ=�8�L�q�z�X�(J�"�;�'�����a�]:k�+��k��������y��e�v�����U�|��ۮL��$e�ͨ(��6��Aߔw�?�l�&��A�6���E)/2�-�}X(�Pr�{f���r]v�e�{�8A��)Ц�1�>K� ��Һ3�?+�J'Xe|��k�?Q^ˈ�{	�P�gV�1���I�3��?�ǚ��ɋ�,��p"�GW�I	Y��\R�/�e]$]9%���T����~*m�0��-�EL��W��/0���.����2��f�$�3��U6��w�"�]+i5I0�tO�nP!�F�=���Rv�oS_!�lW|�zS��<�9�Wn�)[k�C���Lf,�@�6���%n�ϵk�/��*:l\{�RN��U^h���a!����<)�:R�.�>�s�p��Kϥ|�S��N��CD��!VP\»x�	~��>	��I rl��\TN�ZL��'�ۙO�]��Q_���:�:�H��rC�s~ �ǀ&"|.p�t�ە�����JߔJ��<z�r]����嗈9�����ɱ6=�f9UBv�{6+��& jj"��o3��E����.�����3����ݶXwA�e��"���0���r#�Q_ e��Lp��{�w�fPZ[��|��L{t��_�h5��9�mF(�	�*���I�}�&.#��WC��y�<�}��ҫ6�����q�b� ng����2�,��#������ ?��	pϓG]q6�X>���[�BJL8���We��E�+[T���#
�#���{e3�47�ı�~���&]�'F�D����I�,Z! �HEfV�f�f��^��
3#�����&��L�G��M���Fi)E��rSo��YZEr1��ȣĤ!upWe�w%�r	G��Խ60$ԣ
��i�����G�ٶu f��د���|`91�k� �Ex�$�n��Ba� ��$ݓ�����-�MoM����\g�;�О.%���liw�X�ޘPf͘��n!��')�#�!dF���{��۝�m��5A(�gկB(�*�א����9V��0���?�0/F�
���-x��$� ���O����*��![��U͓�8��V?r�R��zI�Y���>y�`:E�V�I���jH4O�(	��T���nΨm�D��+og^<�����fD��s�5ܵ�u��� �=m5/ĕ��ym���7W=f$JL�'|�U&U2S<���j�<Qtݷ��}5!�#;l�;�G�^�Y�I(y�^b��b̮ax?�'�%�	Cr�Ep:���d��!��������*�Y�=���u��&�Z	�F��I�P8�-��,~������l���9���$�>[�R�$�m�&l�s�8�����e>4�T��	�[�0x�݌�@g)�r�$P ²�,��4Ҝ�I�Q����������{��ګ���/�����^Q	-D�>*�]?�H��:ûY���=�8��A6�\���-��B���$�3>��*'_%�&ځk�HZ?�F�!��\?��M\��v�'b� ��P������\C&x�C5F�E9b���R��Ls�E��,��
&"BL��k�(��~��"|��c$>W�f�m'ޜ��`,���P�k��������I���1��G���J�������� Z�?]�|�X�5f�<�E��q>8��.�D؅��dĐ���i#�
�FJG�պ���Ƃ��B��Y0P}��>uf@j)I�چo����7	���t8�����ؚU�f�k�Y������&RB���xm�ٮ��2��=/^�Y���ie��R�8�z���ʄv%����&�|�R�{(D zij8�zǟ8�.�&��n�["�Hŀd��1"�ޭ�����}^g���û�N�8�%!���8'�:�1l���������\V��o����}z5�I�Ҭ'�z7�l"I�م��/�Er��"Hh��h
ݧ;���$��<^�ԯ]��YI!v55����=�q	�T ����{��<!6i����t��/>K�c��I�W��[��6�d����,ڣ��T�����;��bo�C����1�ӈ�5.K-W>OB(��Y�_8�)z.Z��P�#%*��(�0�����X��Y3A���M�,���+�)�9��\��O*
'�RW��[�%��
���|��z��Y}-��|�&D	�:��ԝ��P������㤀��-���j����ٱlC9�f�&^[�P�}9܏A@1�7ւ�<0]����O��m4{�U��륿����t�xpzX;P=�wG�.Ӧ�}-s�`������|gz[�t:����c��]:�@l��*]4U� ���&㠌��=��{s)BHs��f4��ѩ1��`m�ԑ.����5
hS�z�,��m�'���2ڦ�,)(	�)B'ɎH�0���¯G���0|I�l��5�R�X�ʅ7KFm�	����9�a��{�j�S��$⅋�N�6�Y������h���㫻q�������T��Z���0��E���L����
�G�*1� ��#�uX��1�k^��e�
T/̸K1c����Z����yʪs�c�6�KR�g��im޻����Yi�6�����Fڞ�<Hg�8�d��)ql��ќg�O�#�bed$�"���`ݧQ�O���#�2O��������'��N�����ї��4��y���琣;6棶��	'��8l�ƀEw�{�j��v�{)�߹_���-�.�̫
��),�����f?�_�=(���u�b4Q~!��6_6L�������oI�
����Bau��%©�(�B$|c�vN�j�ӱb�q�1��$L3������������e���wd�t�d��vB�>LӠ(�$!	�`����Ź|�W֡����"�����&���~pW�ʖx"�N����$zϣ?�裲(��=^/��~J ���q���.���-�(vh���=�5�ʦ�Q��ֿ�}�!C@�V=M0���XO��oB��+�����T*��"m�}�p�k6*�*/�cNʒ��U��ӳ��������;lM����BE������<P8G�0�����I;*�H,R�
]���0���V�r~pO-�x;�;�p_��
���ͳ�rtD%y�������6�\��_p��Öqz�( ��ޝ4��4��o�X0ϲҺ�Y,��9��U˴ϩʽ��݉׀4Y��{�L��Q~k�����vT�a�d��!e�X�����*�I鿠\�f1R����즲;���&�3RUĎ�:��?�J��U�5�n�E!�@A�;V��]`#�~��f�19*�l}���^�R�a��ꆧL?�E�a�^��|r�zX�YJ��kc��9�����?R6e�VdtF�����*C!�l����NQ���0=�!�	��kȦ����#�����~"����k8�;���ٞR�FF5o�4���$�pW�żI�&	��H[ fs$f�=P���2#���h�N�*��*j]�.E�Z'0w}��I<Wu
��U��(U�錍�����0�uPb���Gו��d��Ew��@���A�5]�Hb��g��@j��t�F�S����Q�F*e�ur�Q��B�����xXJ�Uh�1b)�O8jVKB�" `��z��k���"�<}�rTj���
�.�Ƚ��������w����m���ߧa��7��FPEW@�l�%Ѳ'�˜�ݲ���PA�wy��5�|�d��e�!|"aOb�j�N?@w�5�@g`��uR,���B��?J\*GG4%�)1!�~������p� ��ې�@��.��)�)z�@v���f�����.��܆��w>�xi1wg�h\�u�G��`��ɘ>O�e�DԘӁ=�-yGQ�f��(ƃ�=�Y�̰b�qҬʒ/�D�O��V�aꓐ(��1���> Ú���>��Q���[@�&5���H�v
][<3�$��_��oWR��Z�J`M[n0�͜�F�5�n� �n���/������)`3�����;�S9���҅�O�>>�­;�}�����ں��<�cB����f;6�4�|'8w���ZZ.̋Ls���|��]���yu���|d��N%d�V��@�ߍ��:��^��1\1sW���u/,��o\�����C�aYʀ�i+�{ tt�)�"��7Z��ü_�6���zF�">1PAS��kO�N���p�0q�-Oo/��P��m`)����ͼ��8��}�E�>T�c'I�~o�=|���-���ʦb5��!L�ͽ5�� �-NG�;��������1V

Jߒ0�&#=��	�Dc�X���+�T-��+�����a]�)W&XRjF��"U���D�Ұ�hgŤ���t�'X9�מr�T'������ܜk��t�:���hR˙�b}��/�
'���hё�o�(�˃���'�}��}�o( ~���)�����q�O	�팱�ٛ̓��Y�$(�S`���`/R��y_�)��?=ޅY�˒@^v�.3I�RDr�U�����*��M���9�?s&f���gEl������=��7�C#="G�jv�����Rs*�X��Y�6Z�|7la��$m7V�G]��1W:rE�meg0��!0����n`�t��^=ݽ))Y2��[�3bV�o�h_	�m�d1tG��S�#G�Dymip������ֺ�
d��5R��]�9��Ÿ�6����iV�Z�al�ۘ��}Kp�������j��?>�%_�	�n�����a0��G�nX/TI����Ehd�m~ �����_x��r���s�f���ڑ��B8����,$�#�:��v'}|mXj�}t�������$;1�4��&�ډ��{A�O�V�s�s��AV63W��JjڇC��'K�b$��#4��o��Z��z�d<gd�t_��\2��v����Q����S�	V�)��L/�0�h�j�r6���U@�(k�"���j�������m�����(G1�0��(��D}�{��7:9�p3���l��0�4�#~X!�wLt,E�)=�����s��l��Wh@��N�H�=��/YN<�2�_jo�6.:��O�)���w���B>0٧�( �o�1�� �P�}�禧W�I�%�-0o��(Y����?��K�A9}*S�p���,=4��X��R�C�����0dV�N~g�IZ��!���_��s4�����^�=���Viw��r��uB�������{D,��R^�����自+��ʐݿ�P�(�A�t��_���+Yw�ʹN��83;�o2>���^�K`��F*�Y5��TB̈t�6k�Z�A,���'#�/�Ӹ��K׿E�[!���_>v�,�p���thdlɵ���+��j�*1�%��L���7�P2���)9�&�W��g��������i8��I�{KL]O�aa�8�7لN�<�`0f����@��h���@�T���̷5~�?���X�s�m5�	-�EA���d��tt�,�y7�@ $g���MkF�{����3y���ꍭ�m��U�]�Ό���/I����Zjl�,��]��� +t���Y��*A�l�j��4�m�D�§5����Ю�e_�~����5�ি�e����M��C��=I��{I�)*y�6�iP�����ϙ
G�����/*� �.�s��/� D��u-��)�1�J!�Ia�P�hz�����)��	��xa���Y�¸� Z��	`ϩ/�v8��MD���O����'q%t�Nx/]4�����4���dQ< ��E����,�r��s���v��ϯX8M�p�y�j��Ġ��Gp;I���c�s�.|Z%^�I�Y�������� �Bф
}1��k����1.��hG������9���"�C�k��?1�TA�Y;lg��vY�9��HJ�%��r� ��$Q@��k�{.��&s��Fcd�GT��Y�^!v�����u�7��t�K�ے#�V����|�k�xZ߸vV�m�/�mS��ss�L���������)W�~kT0����\w)�|P��,����E�?�9��V��B�+4A�ǅ��ۦU�"�(J��6fB�D�e��p$&��Ѥ~˰#��(��1�83�-��Ȝ�@��A���MtW��K��X%�������D�L:�c��'�]���䲀`��/���D��M����'Y?�ol�����
���{V>=�ۥ��=�o��9�oPE5�1���u`�/Zۈ�h_����#Zߧ�<cg��N�ej#�!b\����#������rӪ�v-+yp�5��Ы�'o�L *T��𵘍��-}+�����w^s��@#�P���s�`J�Vl�#������߇�SW���>�E�/%;o�{�^�Lԯ9�~��#��gƂ��?��JDa�6@���;D�����2f�^��,�?��~A��J�Hdi�(�"�R��������	~H�;u�2_�� 5(Q���M�ֵE:�����q9��^�����A);�mF}�F�oIV�o2 q��e���O�ǿ�� �����(}Ȧ���2��)L�8Bd�Tl�"$����^��n︩�}S���R{��� �E��H!�2[5o�gmk�ꍇ[T�Fӆr��hM[l`�':=3 l���7p�<��ߙ.6a�JgI��f��C�I�g�z�.�L�Fݻ����C)gi�s!�=oS�N�z�փw<�tx;�&�̡���g:�)��T�� B~�R�F�y$�Um�'4Wm���?6q��J�;o�C�pL�
R6x�8�>HsY ���HX��{;7ӜU�մrg��$�,�<�?e��5��>_o�*�,a���g ���G�]kmP|H�������t��BV6�?<E�n�BUIًA������������:�y(M��QKM����2)Q����l�B�jU<{�����7&G-4D��<D�:�:#�-#�K��A0�@,s�l��U�-������>0P���-�b�Ɔ_����l:yWD���ȿ�;j^�M5p5t���qA��8�����s
_����N�k8�%h3D����Cɿ�c���NQ��TօfI�֚�j�&z/+gr}b����o�����ڞR�!��	ĭ��.�M���-o�a%Io�n��_��z^��m�%�⹃��_����k /ة+;U�&7�TT��\��m|�[D	���4~m;iQ�b>3듫cD�%b��LWAi��<�xd�� z�{��>.����e���ױl>��ز�o��
�s�؊	5c�ӱ�.@L��@���4{W�CدJ0d#��"�Λ
�}C陒_�&]���=Xv�!�����jͿ0�r6�ph�
 ~�=��d;w��fL��ي/�9<��g��g��j�%<غ��4����(T�\�
��ް�E��5g8�6�8���O\v/�8�HhO��N�� Kצi�T�S��~�^ ��!� ��$u�0;���.��1j��c�܁aʺ��ŧ�UW�Od�<yΔ��Ab7��������H�g�.i[���s�4��d1�����CŐ�F��UVV|�:H����U#!H�{�P�����2a)�]ި����j�/@��Ha�ߩ�T�r��h��}]�B8�h�|ѯ=D�Y:�>a7�9��a;�S��g=������i4σ^I\B5�tls��j��
�&�i�`��$�<���׿�A?�Da��p��lr(v�T|����Vs(*О�C�(��&�b�c�N��q:��:~��?u�-��l��x���M�0�����`��+���Wr�PY��{{��k���9F�gv!\�����m-<qq[�K�--���V�{��r"�,�������=BP�A3���|l���<���R}*Ȓǂ%��^*���+pN���F��tt3��6��F���Ǣ�*��_��C&\r�ceu�UZA�@���&�r���{y����LvS�Wϸ��"�GzL$h�E�J��u	����E����C�Yӓ�D��c<��Z�L�Y|*쇊x�8���:��C�����86�̒��c�!����M�Nm{����*��'�4-����~}*|�K��E��5V]>c���ȭi��U�e�,�7E2}0G7uJ�$eS�,��{��S�v�K�Zq���M�̕.���^7�k�<�\�;}�k�Ŕҙ�n�����'�X�� b��M<a��]6E?w�zҚ,i�����e���X��x��n�Hq�3�Hi�{&ҎG9SRL�̤���{�2����|�A��=�B-'��j�p�L%-��R�_+��"_˲{lw)�W�/�gڶ9��gh�>R�(3i�z���!�V;8S���|?�Ƚ��J��7;��bX�_
����I����nR$HIR�Z �v�����ė�i$��}�d��MW�Q��b�=�9E"�(�����]��"�N�`e�1���`$��I�yj5e�b�Jf}KЧ�m�v�"G�  ��zk�d��햃���Wޛ�d7h���m�x����s�%�ֿ�vLu�MF�0>�x_�mK֛�&��ˈ��91~A&�c�\�'�b�p�7� �hl�p��r���35B��� TUc�SVP�xu'���F�J�ey�O�K��Z�û�8�? ��x�t�%�rZkb�9��os����֖����k��=t$L;��K��k�g-�.`��Y����JT�J���! �\��4NhR%���.�
�o�v)�7�
>4J3y�RD��r��DC��6�@�~�<]hh��N�YmA�A�w�`| 