-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
09GSrOLoTOAfrc3XaFy5Iaplwn/t/hHgtsiBtd+1affG1LAfORid41q4214zK8RRi/9F1RCAFeL9
noFy+eThP4/HAjCL3ODNGEmqpJzXJkOZFTqkGVEPlIGJ4rzCEUHcxz0m58LqcfqTgQwzPg4aFTh0
Joc+9VVGtc/HnupIgwKblgIWT142WgsQD9aCl+RQSX6pkZUQnFIURM0yrql7hg4tZyLMrNcN+dQN
PzC0+fm7Zq8UiUE/QmMWjxgPkRPgqZL7D1kT+aJSI/2sqFD/C2f60Ru6VG5pMeXW0B2rGANJU5AU
w4eLGQSs+VurEBX1Y4pAN4NQUQc9hpqF7dILLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
HHcW1F/qkyZFGpVdqoF1WtChF+grxD7VNHm4fkxnFz2I3gMMO121+47zGHkIBLeC3yr2yGfO28pw
7Cx5PEzPFEP1DNoa4nXqL84WmnU0nmKbspFPjbq6WsH7apph0NGnDwKh1/MNwgnZmIbt4IA09YSd
4ltW9lHO+2Zr1FRu3QyXWG0hJkUAqVjwTDojRyYJ8Lmkv1ZOc4tRb595yYbyJDW9q1Fhie3Reep7
jp0fEr5LA3likrHOipJVbt8tf5DnZq6PbD6K2ZvfpeB+ZaaE8AFd/vNaIKkIroBv0oyzodtCeQD2
8SnXst9MYrlr28MHWF5TNCa7fYgKpRgYE5e+rfo6IUQF9+wa/LoryYKa8KrEB5yLiuW5sQB2UFrI
ckLZSM34JlcRwbkrb/mf8SgaDIYF9brt39tjVnHDKVsa6O66kF5MqkbjdzOd/e/tyYiogjF6GMHD
SGpNvfYD0pol9Zmk+o0rklIaWjQfv0n1IIbciW17DY/4LM19rgr0CekdOX2QX2H1Juad8U5yU321
NKABf74azJNdRQ228LINEon7mRdRjM5iJ6AWUOvLOpOYJU4zcbS3f0w7O5HC66mG04ucgN+e9/JQ
tn/7dm4A+j0KMKaYR3jAQKU2W3Ui/m7Sf47vJCeTKOmrWQZUgzIe0PNM778MRWGfl2NHmZ08RZT1
8p6khE9+fYy+sWRbUaq8wD6AjXxc5yuRj4ChWISThUGNvFpd70etOaqAFZlO85r+L5BIsPd60aAZ
E5A5ETlxHRKe/DUDWoJ6eqVLQruTAMz5wPuQZXhg4gNvCM6C/JWmr8EfpPagIsjvk2890/ssbwdS
zy1S7Ty/i7ePwvh+w2NNE4QIywU17LKunriPjn7R9EpoRTSjwTuLYxVq6vng0C0IuD9JLnlfRATl
OjX3nMt0Zzz4x3M8fl3jMbr1R8cBQxaJowmiHJF6mzbpEt3CTXFY0E87md08HKdpTXsNOEArPvId
w+nfdd4TDBZEQEVtyOQXmoxJGf08UkqgrOvL0uPSXhfxmTCTrh4JF4c6QISA7Bv4ahHMPHhxCPF+
JJNQyUJZtgHJ1B4JMFBwhFxKGN+NXGnzD0DbQhh6UJc3CnAhU7CsmBujl2LqGQSXX/wMER7zKphN
ypnKzOIgY4aJvFMxgsT0aISynheniHAdxA8aR2tQb3/VFJBWoHAMb0GNPe6Vh5XwXcB+aJrf/kXs
0ozfIP8LdQVsfVHG+bsaY8oSqvzyz3TP7PfcTK9k9zPMKaB7b8bKMDHFe9omOXOt3Ivbmh7hokeK
8na17Zed+/mmh8x5l/KXN2p4jVZPykDPZ8bnLoONSA6jG3YzvsZeMfS1twVXHoF4dUQctWORQ1Fa
bCGYYIHpjdwPq34ST0Bg80aNnv5tVaij5sp9/Ns3Z0+/RNVAU9caP3Y7yociEQ+/2xeuj81LZoXq
4Q4E4qvk973MTs6+EMwqR0Ap/Zkbgxcp0Y/vBWzC0IclnNriXYu41LpT8u5FiFpIAY892/NO/BRD
CbeKuCK0P2izvcWnBJQAfwEOTl0c4BoLs7AATW59jpARJ0myHGrxHWVQDgRle/1kjtcnG/HbJ25P
pDAFLiHOQMDmyUSMOIpmyf8uxLhVeP84qBVOJ8CvCJ/DH2uM7RoVfIL6aJqBW+1TmGDj9q0A9X9o
3dK3RBs2dKb+v50UrkJKbcnIvyrhWOG3BGwIMyMO3hweGywVLDsBBlaiNYONWjQT2A7DW8OQkiKp
gq5nMxXVlZmebpvPp7s8EX7+S6V0LNyt1/hEj00miOkzMgHqm6ms3uPUNypipUKrpC+mTrx29iRd
TreE8rEP4E2+0YmXMcM8yALLOhLtCl96bV0ROcS6UxLtjJExC2XnBllxNgje40mFlh9ewltSXaxj
cY+8gjXN0mdOyYgxvxir9C+FxQO4yLY4MsBtYV1c1DhPtCONkqIly6ITzHwV6fiPxlTUqozpoKGG
BqXqKvz8JURsaWbTKRi0Q+CtgKJC0516ETv8H1nI8YITbolmqt55hdy1OgckZ99ZhCq4lOk14I/X
ZnyxVMQehrJX5btMD9773O9GARJJkC5ZRKZNnfWi3yElycjUWDSuaBCoGEEl4+K0TKL0S0xoj6GQ
XJfu0Pg9qPBapR0rmFyJ18N0FZBma/VNcJbOFe5FCCB8AIFMB+mSoaQlDUs1+qggu/uI8uBXjTd7
KV9CDeHqK9fwAXw+HVSiXEZHCbzmw9/RWds/iFbwUNzTpJ+YpDn4hvzLanXBI+vVcmFN1L5yvWyK
PBff3wInEE7u1qdtisWvNrdBKBhwwmWlVRKvNz1CVR9LrMl+zRyXm7jzsCx3zwF/OQiMMjiR3a/d
LLRyMp6sbDlj4d4KvjASbzLjei5Fu6/nyB6Q0AK39DsmYb4b6DS1EYfwugv7I3FEj4kG6SvdxYQ/
gZcpYm0KNVApNDjfb2JZmCWf++NSdvdveBuNN/FVCYkobAlaEUE0VZmNjvtqPzhX0wIM28r0QlwN
maHfXCxfV8AVd9axSxQ3IS0rJUOawmvl/eZekCrrwKQEUnxJLgEK98yZSJLq576Ry1wE2uNNbgFY
+7K1h1n1Bx3apn0Jv3lOltzZ3aU2/naso4cVgYKg3qdq2AUalnaIfAZWrL7W7l7d5tz35kk0vNgx
7tq6PTD4MearHjq9phTANSiE3Tn8x5g+f9pv/BbHvekuNGhTQoHNdsm37VUikbBStGSeFQ9Cjq2G
P9tcjU5+q5knFRJnBHlGawtYDwe8QRZiT0id2alk82VSE+SZ2t40g9rkk7Uvo8Z4F/8IlnUn+sUq
NErwzQ4zukfWKPlEc4ylSNtcsFeSYCXlLtRCS7o25UAuqnGsL+iwORBIukYhny7+fY46THZSDWGC
GLz86pKFivWNk1GI9ikO1gnkc352++spjd/TVvZwhg+6XBvY68ai/eKHtUIxGMJ7SZkNu36FP9DV
2z8flOjerAuGAgc/fYgQ1ztqpDKO4FyZ11e6n6zc5cpBSGrReSKrUAtGU9L9gaNszP0GDIvwickN
xKNikrR3/Uyw/jUmu6pw89xyBPTsgx9mvEVPHZLQinhChanhYsxbTKS558C2HI+SyEBou8P5J/F5
yFEVKwxyf6+xXGBb5AVfoe6EAyUJubnO1PBe3CqxAvZKBwT9Vx5QKGyc5aN14UXbEb8qH75b93b5
7VkicgBuFzdr8Zkmm9BmuR0lN+j1HmQggTvm+HmQ7FTMI2ZOPxdz5T664hpUq0Ff4ItDVu+vo28O
u3OFyeHiTblFg6YUZJFVO3MCfxN1NI5x7QsVLWrr8k89x5/SnHVUINeliNtt+OwFx7QJU97W8Yuh
qhN1Dzn3aNZwYjepPkPHnwqodJAmEGgjaj1b0VrrdehCfIqKq531XoZBiXf4ivWjF21+aJcb6BNN
RGTtCb8o8utNrqt0NQF9FmkRMki/wpmKOqZ0SbR7ngwVxu+v4v9LiJCdkOGfXwbfMdMbOwCqLnOC
ORs7pS7xvglSu7Df8s3f+zvamcHMzwleupxzQTCFvOXbqRslP4JAVm7U1EUo62AoDTQ8ZVloIugh
563ZOjzNU51L/KXRkIt7ZLhO2IBam9is53bCXeRB8FrnrvTt4bidyVu9K1vkf8g4Ru92onQXXzOt
kyUNFmiXBQElz22FhdA74+7iDEqMjRVl6kO988L3ojp25nPUECuoQG8E/Qf5e2U67OSM9C/sm849
LYX+FFZ20qbT7oOFcEhDwRyne2y8D70Y6n0/jJ0TohU8ykP0nz8bVZbIu+CWfrs7SjgmK4s99PA0
bRH7XfTqfUwxdZJLJdtBDuN6Ofx2MA+FRlJaCPfFb6/IS++4SnVsQ1OEysI0K28se0ClPogS2edL
qxoCzuhA7ZTOGFP2sN0zTcr0HkY7m0OzpsGm6cx5Aa7R97X+qhT/aN+iPMLPrAJhE91TmErQY3n6
yF67bro7t0SYnx3b9RiEbBRWhuc9MeTFSihELUKmihWKTH9wexrH4yTkvFV7a7bfNl+ZYvz+GCTr
cE8wPMRhaXg2+/sWGwYUWd8juoyvdZxklgeK5/ISiorclvIWJDlHAdvyAN3awSCg7hSc9TRJhggQ
UYGbVbcqRsgswE0rTRwrL3Ncieanns28XHMgR4mSs5Si2zXz5/8yJlywsiOqOiopOi54JlcEhqSw
W3PzvHiWWx4mmaX6P3gJ0HKsFZwI8txD8MECVt+b2gK6xDRZJZvREWJNOlZNfqhF4Btae67+w1pr
zx2Qtnq3E0O0x7EGL41iwlAa585NtwaFtZvnUBqtYpYD/lUi0qMUA6LCjoqir3u5bzHA9p+nWZ6H
xRWs3nKEKt6NN992NxLxBqz5JTJTK/Bjd+PbwAli6YsOQPyFOy0pppL6gBiMgtdEa8Ax6rDKBF6B
z1Cs4B8KHs31Iu4Yf+ViGWL4BdIZcAmAbOwJnHFAwdRn8VaK/nul4Oe0stwnohMX4u70mxxkVQbD
LLbasqFiur9rycHyFtr/9snmvxKuuF6WQsL1FL5frq7TWphoosNnu/Lj7Tw511xVBvdTJeuBPr/H
hQ4Imm3DyVk1oIwTVI8m8i0jNgY3MaElqIasoXTnBm6G+0V2MIpLBDAZOvLLjGQZeRHMcZz7Bo8y
aTmlFJ1m2Kw8q+EtdmjtP2dWhnx6/d89ZOBJF87l+nme4E7+0CAPuyg6kySGUWQPtD8FUu9OeEvG
OdzKiKYvYARPA/mtwWiiXtu1rawt6UsWUAwY1Zr8z/gtEbm2u75n/62O6zs1ETAJjA3aZywp5npP
ehP2TJIEzN3Zo+cNIuY6o7Hv6jtnERxAg/IDc7FKNhBcbxP4x6+0PeKrTlYFlIS6qTwA1C9iwTAL
yxzjrXSzr3hJTI0IMXpyzRKYFiDsbLLSEli7424pSnULtP/5MbY7GakAgkzd42sXwwXhUfZVCbus
kUYSC7kNxHvwZ1KCpsEH03uHqzEQV0Aghtl8DGrhAp7pcdG6ZVr/W4Q8WSgYBH9T6Zm+ZRlAM3wt
0GbZMgT8jLToM7auIMD37pigcWvrI8LU4tlS402kEmjvG0o0Imm5z2NKCPs448CqfVIutYW+GLlZ
mkCBy8PZpmBjFmmcvhdX/mZ8KcWNGnIl4y4CU6vxUs6kOnCX8v0F/8580Lrmv/ttTivk9r5DYFCi
v6x+eHxN4zzr/0DlQjrYw/65dm3gTGSjhUuxs07wNyqaPAXTOYBTgDgT3MvQdDC0f0MRuAHm98Ef
6gxjIJxWVvn2dhdCaazT4SAlJUeOMri8ioqSXcoiPSalHX3ame2bTq7dlvGZem8y0ayUjwgkqwtr
hCQwhE66fbdNQkyAeIMB9rPPgd+9m1xUi1IVzWLgOENUzvTPBALPCvXT4tGgn3xo8qxbdFi0D+9I
bDz5xo34GodMBQ8mvgHlzknjawEGnrcrRY7HFPw45Bn9IhkWaT53yJrWLtuvCZvbhFLrdsHHusOB
BJvqGhwdCtsDTwjXFuxx/La1SYmGzdWH9aytTgiT/ML2ufhBD6Xm6CmiBsunsHeYeVwlDCF5WxiU
1TVCZ/dGE2zSC53ps+J+PgswiLHw17hYLa2Ts/7RnIaJE2Jz7BDiQmkaWUW9URqr8OGwsVIeHhf3
rvP8HSRy/L39EqvFefYK4oATuTRT4PE6irHuXxO6oEtFJVaj/JGeWexcc1+1jZX8nmQ8rGmWtssa
lC/NnEmpfLF9ndw7MP8RVgaSPo4zS9wPrrm/+qWyd7eCOdb+baoPgiqY3Pve2T+XCGAfwTFmkDGA
PoOJfhfBW+mkPVPAq9x9nA+WvitIea2sGYDH3cvcfyudztD5pAjiwbMWee51DYaZGvW6HizuR7XY
Oc4BYeTdEM9l32KaxDvRMUaIIBdlT/YI/lATzKhtxrjdRcG+T9X4UJOUiBrDfhDk20rBgT8TJHTD
6b0Np2Kdef8Bg13ZlwQSUMSkuZq1uDij1wdeo5xGc5M+xv1f1L2UCyLXaziQfeyelLJl8Oa8XJDL
fr7Vb2hzapNJGPJVuX+np3H81fDYMJLAK1lPbI5skER5G/PlKFxGTsLZaig99cRlvRRZ0jgo6Wnh
6jKBG2uK/VvLovqVplzVv0Uswo4B57wQJUbm0jJNVi0HVf5k8p/lmWtJxK58sXSgIFP+qZKz5BOz
GyNRgh4k8T4dZuxn7eoqRaeXf/YMb9+pnKzhXn0hMDLAhcKPDpPlp66xMXPm72gwC5Xn31QvMda8
QeRm+S9fRX2PCN2oUIF4ed1e8WpepfV+8NJGK+F8qHKq60cMDdzrZ+2h7+lCJt98xTUpqGXKTMbG
7RpDCzeH1E+rMUsUqnibRwtEB2W/8HO+bBN0CYoLQLy+yLD06peWeV9LlKlORlLvvB2G/2XMKlNb
xUVX9svWQJGk80vDKOq6hPHRO12B4ZID0siXnA==
`protect end_protected
