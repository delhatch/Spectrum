-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RqVi3hJIhJXUtCsuh+JhCJCA+1lJjtweqDps3MHLhBFTetXTE7J277yUvSEbydOEUDwP4VS8uWSx
dy2ERKy0gE5B8qhr0VKxr/eO9JpbOtT2FydE4f4J/UN7pF7q/DjDQPQATK5fM2uYPfDhOyXcF/bp
yhD/g+aH98FSF3/b+NqIDgonxocTV00HEiZWtpcFsyigRdXp/c1T1SXFK5xW10v8f5XppJ3arbCD
AIeWOLvMGNCz5EMPiaL4JOqA30CPsvrJkSyhahROR8KL27ehimhbKps2x73nwkKKUze+de7pemKl
HXDMpESLwPxqIt6ZQmSf6IGjgCjrw/ErIF9/pA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
w+RlST3mVBRpaTdtOuJD/Q5aKn23P3IcNz5m0Dxkebb3hQWYw4N/Q4Kmt3xgICmBq5gxVZ5iTuYY
8fZMkzHz8PTir2FTPKmdjAFusTqwyPQ6B6wXXfMSbHAii+hG/PHYrBGFlWUgLMdBXgoPq69iIG1C
fzcFli29cyRrb/ibMYantR7P5szaE784YQF8VmdYYxduxab5zkqaI667YxCGYgPAqGSYr5JM4QpN
aP7yiksoSFx0OUBsTFlCXeVTRHIB8w0HgM3oTBuTDW8arWL9SVhyiJR2NNSG4HF9boXWjYxtDs04
5B1zX3DiSbKQqayaXd5Z9/csDB2rDIVTWrdTKQRRqGyqkqCzbAnPwsT1Cf1ES7YAFFvM2xZKc631
EqUjyfjee+Gj1ou6hMHqmRkzx0C5S+d9Pog9iTRzFYPm7SS+Z80zcyT0kP3+POfysXHJMEhGbSdB
dlr9/l6rg+4W4b9mXjbMDtnnzpTgxfBvMN+Lht+yk301HZaDYhukztZYG/3rc0cc1HyXTFdqzQso
VL8HyOHv30epy3NOtbz7w27VuqdG8KIBL5k+ICx4V0KqKCjeHMHK6lS/8fpPqf+nRncdGzDr0xsS
ePpdLWJnWdZx2I7SQuEN6AVeBMun0Ew8edDmjf4jf57QQXtLkLdcSZjcgby+RkP6Mu75Qmx1atGv
3XY/A47PYcbgaCjnrD9Y2vLk2tAgIhIzrKCuy7QkFfLjEW8JlxYVumlRHcx2zf8R83thvx/kOTBy
0ayFymUznH4Cm2hhnsL/oRp1s0Fr0A8lVuFFhGeeRc7Rl8QhzaUjXi4NFQR3RAfOAq4kVombtvia
SbqnbV0jR89cu9IOJVYtv/1ysO1bX7PVDBFTKFwKi+6Z7xA6ICRhoGdp61+iksCQW9Rt6o59t1db
bghCRjOHPkvb0lO2Qf3JAhqnveNcznkNL4fLWEgoyhqZzUUbuc3Ynl0KGi9muxyrHBbQ5bs8BTNz
O/cXKL1guNOngqvju+8FX0HEYx7dxxGk61Y2quVmFl8j8sw1y9LbGYHYDmBIpyW9d+WCrN0raLbh
XNF4NHjPN96CM/bW0szmFxLCVixT2fIhN1quN2jYdOnhajT93WXrsmVD0ymW62posPitwElFzs5V
erxbjTEESTx9VdNMUu9QBO9GmqtXW6vLJIbJRpLfKUO0+GMbH4rzrAmEbOu2fsg8Qv1Vdea2GF+W
TubjoJG9A53/YWCz4DnCZdIvNc5WnECWwL013Wec64dKyOzaJCrmXCZuYs81QoGx0n6XttcWDQaC
z3S7SaMfGJskf3iv0R9lEC5hbpVdFIr9KWH3BBqTfbbM265QxTzbdLd2hDtQqyETOCBDNE00zV83
hnLEunm4cuqwFAj+KCi5m9QumPS/nbT6rYuXIkRgPHdvr9I81AEbsS46ezgDOtXI741fLPTyu6DJ
jkaKrc1yQI/Mn86TGlpmRF3rcn7x19AwjfmdUEy1M8JhZRfpWoLDAxXQz5xmdXWIMehlqyYJi8uM
11eqRqsRehcEeA/o7sPHwEhKV5alN5uRIz+pY3KfvwQpEg1bRYnzaOCbvGR9mv3rWqibR5Bu27O5
4BjkFzZLLfIp5y3rYumR9L2xDq6HtMAfIciR7VI8rbvKdmJMEQOlG3l1ij3oq1hKQbp3FX7BEnxZ
V/roLH6pF7z7gVjbV3ZOtiacZX96URoYUy2qaIBABWCHTuGYQ+r7ntdHuHVpxm9t+gSLe0M/KAlK
Je/QgUbuf75wosMwgz02Fxm/JFMvQdYASsvKhD5jyZWQPaSPs7jYFqmpOZxlGi9KweAQyo/PtoVk
eQRONibjkEhNVSDXsY56vHWTt7tou9+6Uv61fs+HEOyKsKo1zZnZindBNlbSO3RqkMRWtO52aD2j
oqCELjcpshKnDqBw1k0oWcB0FV6ktNR+szOZNvGOlBUK4PkNCQmsBVA2bdS2a9FoWHmzpJZEt1UO
MGzMUN0DvnNX3jcfMbdYsnoKRaRoT1G6MTsR3miHzVVYvT5xrFYfVW1xTaW7GLEqp3VWLp+ZpIF0
7dJnJutUPeL8WmEnljVSlJRX46YX2OgeUfPvQyEZ+Apduap/3XJ7Uq5Qm0WBB/FXS0wNpHgMLzNu
X/C7y/A5janD9q8PkVpuXBxAxPCkvWR3FHq9eD70jlnuHlU0Nms1lGZjY0gUrQO3qVSZZBTbBYMx
LIJBByT9dtJA7+sVhLQ9Vt8P5prQNRCg21tDfrOtwH/RSG+fDzistDrd2494EPTqO4m+pKvLuW7+
6g1sNwhrWr8X1W96zEwk2/DI4HGd1EkSoiYOPx5EEO8tDck3UJyQU5Pht6D8iUEwdP2huWzps8H4
DGY21dqLHxFJXr7Ply226D8uOM5maMBUydjSlUbpbSoUggqkQJ8IHCOPWJlv7Fr80Hv3lYhDCCru
G61VglGmCxk6ObX2/Qih0DBkAU48A3F53NTkxRBaDvUNsEacOgOLBMDa7c9BE2Qet75cKbLBx/Hx
iJQ4qGJ06af4Y96StiiTb3F0TpqQT3/yoP2OrceKPdEKyr+/sj4zQvzsmGQwKRDWGquSCKvIeDdh
KJUMelDsrDTD9ECPYn+Ey7USoJT/Q3F13bBPc3hXYUNgi4COTZDJjsqOVCc5K9Lrvtjqp++DbkzH
DdjHt1KJgQKbhgqvoQNmvqakk+gz3HLC1GjF8ZRxAtiCZaU+ZaZiN5jD5nC+MNknN0lZ+5tj+HVv
0s5HwA585+PGe9PiWhc/pV1TfhZOAo1ZNT5qwqDGAzH/lbfQ2E94zz6wa0fmWbNOloYuueZnVqHt
RBVxxiLWiqssdLg3Tap+/qtIsiWv2JbifMT6aIzf9kNPi2krs3RbzrG+cJJw/IKK+XlAMpVRhKBn
UYhLobXj34m1KeAHVmZAQewfv9LPYB1Q/fIlC7ILktyGbpf3D1RfLnh2Akq9EOtwzeagNKZ5+Rvd
BJDYAz83K1un0/qxT+HXdIR2v6zf6o3ua00ciSgoHN/JLLmS4760AMgj0sNdF+QtoHPZOHxSZ7gq
gGkJPKrVtxk6v5l8UUXaloTtJinlbmRDBn92FJ145ccyFV2VcaArHh3C0p8xeKquR4lD5Q8WHo/P
Okc8LhQXQgYOkNY0DqO0EI0D6WsX7mAZtAAz3STCrLI5jSQFS/ewZjLVHwCXy5mu22oYMAQoeCN9
qmDOG487C9L6X73CbV9+BPLdOQfh0fEmyLD5X/Ec0L/lEHSWQuwULQGN8WcClywy+al3FWTEfbTK
nhXoJtSHhBTWqaOFZgHU3QnQqXNqhd8CTdQhptt6N5uAHENWiAbrDl39fDc1hEGX2AcnqgKJqx3r
ScnEjR4ETHLOkYAL2/dqW/eQ4lyEAyRrGwiEvH0TGJPX1lTzyDwaZ9aKWxccHAYWk4NBUnCBmrIM
GeHlyNmMX/to+p1q3VwAPnwPQ4crHlsfvVASS060dhwqvqfM/ogAUf57fsXpyUz3yinPQ80+cy/g
8iK3zTviJ/LQtEWoZXe7aVfs6gJ1bp1vvuP5HdyLLtriN2tARzDges4HfKqPb/HvWfzxIFasoiRn
VG4rG4tUUGGaQulMCJhsjPTqcbim2x7mqfqTxynPQQqFPFkPmjlbAq1qhbzlOT9NRg7cayY9C0Oa
hoPN05SvsXkpPB7pS6ZTQQYwI5R5rNldHJ8yFNtWC6i1Nx2Hv5jLpz82luCLaGuC02IIjTmbuCQB
rqQ6/+d9QihUNH3GBgsGmfGdCjdGpbzNA+1OLcXSZqDaI12Ve+CbOkmXXwFLgI5MXU8/uL7MDEa4
lmRvqL1zm8tb28Y6Nog7MDkzS9YbYgSfL8eFrH8Ahe4oh7LBLTGIkO82iCzxFwpeGt1pPS9OPEUT
KDZMhd7hH7tSyZr8MabW3Zjgc0CLefiJ7SuOCKoo0Afcdz3lyjRoLjWjp433gGAirbuU63dsQmTR
oizBOYEYm2jYthJ2yIU7YYAJlUDdEFPmCQknyV5dQJCfNgrCjpyL1+F6Dh3wUd5vPs61hvkUzjqf
ITEZ2H2M9S2zWDm345qur3aHM0/mqIuYCh1epmNiQnDVKbMzNax+6u0VyyYIA3sZmkXdVURuLrpq
pDncRovULN1qotauCtEdfGUaQRsqdMAerknRmXG7cPuHUlLB9O9gmwIaJsEzwdMiTqf8lBZ/w+qA
iKJVF2+kCTieO5uwfCBiVlcaZ97yox+aIb2xjxUqv3zj9v+ThsGmq3wbSxXfwORnR9qKJxaRxLHQ
47raJHFvdkO+FQ5NFBNrk7CgUQMtrD5rSTCOCy8a+Foh41EzaSZdILyxsDivTy/Z1aLy3UEshfdP
bsd9ImKWIQWelwPdkfsdeKdEWBZX14jZdQO2UdZRsvCt60Pqpkqo+kOAFHLaDmAOREJQIwXEJowJ
12DiiOql3qexmZ+4nDNbHosXV8OrOIxz4xohu46I0KI2Evk2HrizoJbqQMxZwSnHxZW/WYKvlgfB
ksMwSvQXFmUPsthPGfUGb7FR9OXMpNL3PpBonuO7bcq5FFm7rDVd6M3kOp0v8oEv8Yai3anfEB70
WFaQaFidn7MfulC6GdmwpnyMhEPvyl9558hsHDyXj1/NUqyU84O+gAZ23D9/8mqATXxYKpSy7QFb
yjShba86AP4BFnmiFUi65MxSpuToqJIOW8ov21cArug//YiatHftZYxd0joWo8lo+7rHmzzEewem
vSfFzEkAxK6JHjS/27pW80726RPCQSiwjgf8DV89YWDFew3qxfRBntbIqBw/sbl1+sKn8Kb7qRm2
XYhu7yKY+hWJUaHyxm8v2rRTTvPqwVrBGTytqKNyivk8H7+iDPY6OWMjVL/DuvleQ8VoXNUzdxvi
nmdp9XZ9LAt5un4egJv6ERXi1hKsFPlEh94KrlAENa6XSPnteIMDWySlAyJ2kcNBR+z2k+ram/Oh
C64TwXLv/OGHug3cv1iYT3pH69/RiFAsZYKkid6btYSwqrNTOAYUdKa8bEhJZ4AZ0FsyOCdrV+ZG
uo96IVmGIisojzS+pkdI7x8eu/R2stswX+eEEho7qDtPKln9QPLe60U9Vz5yPZPwudEjr1n05++U
txj2EQqN2g7gMa/XZ05NIpog/j1o+IM0Dbg5L3KoTolua+xfChdzJOtSOD6EdISK4OawF4pRJkiQ
9cxr84GtTfWRisR0rWKtjiORp2p2phLPxyCb8IsofEPlaMfx8yM/L3S/D+uLAPwEhwW1fu/01xKS
9GnPEROk8yB13VCER8gpB6nj72dXGu0DxyF2aNPuiqjy07746/ZvtU2M6HGiQBa1yA70Lt5Wq+lm
EpmR9R210NJGrkh562jOy4k53NXASwI0rRhwwWSJa/lhsItHijABnP8ySZLlIhee1gr93a5YJVwD
1i4axPR8y0v8F7Nd5SjSdOPnsHsaoQ158Ykimrvx0XxkpEYtbgC691L1ndPScGK7jkJrfzsfJiXm
D5bXcEjRaOfzPD77am7gDLH1EArHhlYr+Dzs3iCnmWB9BRLuDLB4a6v/3GZUYoRrzDRLNiycW+rF
H/HsETkENOd78/dk5yE2BaAZwHiPK6pwIXrafZHhUwFiGq9FWRrPr3Zg7aKe+1C2hpJ1ue3MSEwx
oLiQCGqLs7YXeaYhpaxR1DTo/VxGHFeoLDdgGm9jOqDPuzFGf7xKO+AGohvLxxAMzeqlCSPqksaz
C71OS7BOw2DLWrWY8AwPoM0uu9wvZdFwLqMbgGssM+u6DmlQWhNacyru+REpXwIWUIvlC3IswIYV
UBXSf/Hche2ni3S9nrZxwvG7RKQYeZwIyyemh0HV7Q4LkRyHxXDDs8EBbQE/5KWk6i8qEXuKRaNC
wDPnMpIiLOL97wx3h93bjSCyB/OSutnOU4xnkvMRt/oAOy+S/mMQYYO5a8K8OQQxdL7QxHikZIVz
P99CODA56vj23Yg4CiyskefRAdqtv6L0iuOMkbV9q3M8K3W1pk75SX5mspZvdjcmQ1gtpgstBvW3
gIonoYenPxqNxWe9hhqKnOSOfbCkg1b0uHD15AB8p+E37vY2Ny8GjH5Zo3PoXsDCl060Z+N0FoWk
4bWKVDlTs5wgz0AHYjeorLdMuSdZmjIXXQmG0SCsE6TlYVVgDMFbBxIeaBBElKxsyQcGiHWf5uzm
6NUqkEWawuaLFGOvmqbkWP9iW0qDUgTtiuxPOuMbmm3Vi5WnBKmhXMASAftWUhYsSlE61cVJ+5Jx
HhzSCJTn3toUpiuSTpFb90QGowpmRpmmxR1eW0yoON3uRVY1s6tYbsI3HFmp1o7WfgBLPUkUma+h
P5wssaLhTmFdayQokUUcb7o+Vw/QSfH6h1fzRY2R3PaEwWfC7D4aisyqG4KLALPDnH83X9pUd58Z
+6QZLZ3T2ISS2rV2SZxOp7GWrpRYKUu7cgIMgXcJQwwZpWnv2K3yaM63bMQE567ZbqcyDeWWNJaY
m4lWDAW/fQTzJs6YAwp2V6n88+5/1YPIq7qkzdj09xXjv23eZGhoGv5GQex+FVSMC9IYWQrwEWDf
8OACn/2NrpF/YoEeXTNu0wp79CfcBEI/ntxl0vTgKmD0dOG9iL3qSkPEUoiYUh6XnN5tp9vGCuyO
FBda3N3fiIRvqzyaQpmpz3Clp9fGs6ZDNM55NhjGUFghKMeqk7uqAP0lMUiFByn9d3ttnR74fWlm
McK5PthGf1M2RxTk63R6cC1sQ/+IFWRxAo3bnWIJU7IfybOzYXx78yRY6jboAI9NHkNr60Yu1S5g
6yl6eLonj9O3kdjyIehqbwEZAbm7H9dFuBfM1hFUdjiYqL3EfHFMTTgMD+eUfqsk8XkBvC78w2+7
uRe1umwN356YHsUjJzIdZA8Yu2YcNE90m9QABuEM2kmKHt+i0SDKpQHKJIQexRBeH5G50f4Dq4Yn
qhSf6HePuUNiW0ShXlob6XTnS/eKcSX60wnJMiQpKTUOwbx6kqfSO+n9AL9Y/fZa1Cg+xuGDlFjw
/NuIfJCp44vLEX5RvDwnN/zpcF4nbKmi/3IxYlqT70yPmGi8qhtU/bvpCqS+ydl+X9hIdvQNSRBG
3ZRjMjEANJKtIA8e32FfrTts5q8qujSZ/xaofaW9mdoapwawORt1fPgBbqotm5KngN0SOvHT0csS
zhehYmWoUbfUDNl2EcesdqfWZqQuqJVKnweitsX5XfGeuSPQWDsVlLPbLy7wIN5wKhriaYxrtfYs
CEkbZohnJQOve7yCpkLOSFB2zU2eRQ7SDT0BznhnHzdMpg+6f/oj26owfV2GgRmInNfjaYr3tobs
JG45pxXVBXYdyp81ZbhmnK1Vl4kJ/a399nvnpIBZsPzGxdoY17dHRaXdwfKPTS2gVPMZ4g5SROkR
yHHmF/tTeDveAAOEorYo3lUaCTnMGKvnm20LgVQuqZfUs3G0qZ5aYitujATb0xeYQzySNlYsvDFS
VMHbJ/cti2EyVc8K/GgGetaWM0BL34lY1qxDNzkRu2IyPMZcgknd19nVrGBLiOMvSPS+lHcGdCAX
00Zu3iXqkkuRKK8P7n2lH99Ty/Ra9HP6dDsF4Zd5qEsyvo2lGF3tVYAqH2mh03rgWiJUix4V+37X
HhIMbSrYBN3nIo6yMSU6vnA6WwNCm2XFjtYzRXr1HP4E9+5iGGrakRWjKYNooVBjiDRp/W635Puw
Tk3B9TSLlAfLaEwD5/lQLovWKE3TP43INCwIxrPas9MFJg5DjsLDFjE7vD1gs91bRw5kpxIQHFuZ
JWdZp1UTZzBuY72I8BiYHzs2VFktxNnUnmyn0QYdSeXFO0mC5VO/4fQ8NyGLEvRg2hmvClOhyl5+
fkX+3U2cRCI26W3TiPPtUZS69fpH+1N7Om4kwL+TMK8PVdlQlIlzBesIhGuIQLRsNOeh7jYl2SHL
RoN31r6azJsBDCQZCIJbhTGdJidH/Gfi6BrFCSWylY2g0FGgzyDYvoWo/NnCVKW6cq/jMP8X6gHB
AZvTDI9XKDkcat7iJXEyAuv0uux+L7exveOlcqEDE8ljetZw2AjbYy0OeHAfRslGGbDezDYtBcKF
gwIgs5SmW1g+h8AySg2BDd2ZdVD93vp4E5irXaiGoNYF3AHq3V2pjzW2K+LeAdsuygyHDir6w6dm
GxapZMEEfToKRTwiwqNmdtyakP1z4ajdl5CoT/wOyER8BtsDzzeMyVX5NpAfpxDfjwolRRDPfeFz
TbgUqTj5AipAEjZ7danOaWieIy3YYn9eOqWzklpwGejFKxzguEEwJDqgti+ITzhVyCN0EvWa+nsF
CFPD2p8inNi5q7REc8dxX3ibHiKkSrnTrjp/4aB+dcQYG2+E2FC+SY36XpLHdzFyQdbQLg9STfq5
8BGT7TFtgQ/Bed4DSsVBbsvkr9cUM2rhN5Oic3CYUPPx32ufKl4eB4V0VXZtnwBgnJnGTHxvkyRj
dp6BW3Ewuags0ChjV0USFTyVNOc0udfMCx4A5MqOFDP+GFmXANYJW1R/LIPlsY9RfDFYrsCq7OcW
eps11huFZEIiqyBzdcR6n6kybZKusp1bKf3lOtFW/m9rSWiHF+McuWQZeYiBljSmX8Hcc9bl2iJ0
k+BDO6h72iXr3G/0SFCb9X84eXnnMyKvjGSaciMbH/QDSdNILcNWX7agydrE1gK8YWWtOkT6WPhA
NmjuJpXBhtQuYdkZKS93cEtGOY52kuJE++89xfmumrGbYkcAsKMV1mQ+S7USA9sTrIPoAQbuoUaS
xStAt2Ur8+VHtmx7mqHBBBFyDVStXy86GaGLq+3eOe/v0lToVAomFZLk7QKr+h1TDqqNDgc6BbVZ
1StgTnlo04+Sr1CGuY6OSx9YDi0izZnldg19PmOmS8mj1OgNERDwjaw/RtVAEe2Z8HBBKqtZSoN8
IB4/iK3d/rbtqNZa4wAjhbbE9pTz+gNzpQmThiXRcyGOblGg73MAPiDespXGMgoyqjs3RF3YkJUB
W5U4vJtv0OQWeVzXzD6nGq2dRSpi2/+4rsUugkOGTmJTuXZJ/OzvHbbBHH7xC/jMi8j29lSXivik
wmnf7lARXtckgxLNeyNvp1yRLA5T6pAl04HLl1nBFkqenTsShZQD64n3UeCeW4mnuChoQtyKsEO+
HPgoCSdb6jrCMm7gRfDMhL0vHK1+0x0emZJIfYD2dg7WObigtk66UyF+AqEZicaZ5sSBC/WZCWaV
ITAStGQpvPuyIEj6Mhu0ZpTGLTpnf156xGboDeTzI5RvcDCAT92Hlh7p3XetWC+kkG3hEDsnuQXt
5EwKh87NdACe4Bm1w4hjAja5G36NLbFb/w/dacF/7HjZGv6K9N+9xfjK8QxZ9PGkIHUN8hzxSAoU
5MNEPG+PN31eGHLkZ8jXgxHdeEMIJVUPldQP4l9XwCQuy3t6kEIrCFG1UbbOePwgFSRbCcDb0vpd
rM0AHpxGVQD9CSYGkh5outyCT578gbyp5EogrnqtOGmmNm3yYoAVv2KU0DK4ASBdUFC7rXuaZa+q
VVh35g8QLx+2REQ+XVa7xLWHht2FaeH+8odcNJYT/F9P9D4rN4FDufoo5Edq0XjdtCrOfGRdsmlN
uOAoWqWd6zC2VO4QMOjCs7BRLh7cxIl+g1uDxe3/2DTaQxwFpafEjftaexY3kxUou0LNwOR4qygU
4ekt05YQkaHLIjwlU6eaXW+JfePGyaakIRQ/whaMvQGbe2upWGVeEPKzDumlZiB4PCrQzjNQf32C
cN196E6vZtJ+1EWX5IgG4I7o50eowXZ1YbAyyLWOqw95/7mlqFwzcJAWYyshfqqdufQGqyDQQwIZ
12tonpUMN05O8D2VqBdjXNBB5udeWCrRz7wugBG5W9nHPzrewWM2rg/b1XDV8oTGE/VKe1REinbu
x3fHV74SlsErZxUexWhYCfdAoK4d2xStN5CFiqiAsEUWDWutMaL6Jk0XSm8CWlKHgon0aZyVcXTw
XQNCoJE+/2j2nIsPzIcsJXEeXqEwCQ4jBUW7t2RJeal8Zb53Gu3Zyr4cO6WNn/yBxSs4cNfjgNqi
o2LISJ+NEQhJwpA+smYJ0ODE1aJx+DGF6ULZUlXStm081Jjs9u8ZVXx4fSO3DZ8NYaEs7q+mpomP
WOJZZDPpVIV8lkSGZPTqcBxMnlRYPkMbHnVwVIRSeP+00A2DEcK6WDeQEUYwpw18nW7HgqG+VUdC
r5rjoVTkK46OV7FdZN2TmCw41h+TPlCRms9Sh3Y3QTXDmf7WzhrOjydibpQZRtlQxhJVqL2pP6Oe
ohH21a5GwkgzwN9G3mfRTcWXJBK6ZtJiuMMDoaOXdhSEOHC4YlZwM/EpuDmgqUQr1GkT2QcK965A
jVgqrPMqR3hgXA94LwU1ATYxGYP1xMjbmnpQ4Dj48lUKXg1xlreP/GucU//Paf+5W2gZ552gHilZ
K+7IfoJ/ch6lSi8cQcF4v+WN4LTaWpC5FFQaIfeHq/RfY3yWgg1yYXAnCG9On6QO692E7T4nLnKv
62SIb7JwiTE26MLunPcdxcdp0MvT6kp2iSlnbu/B6VjIfTSNrWZAGm65MmbwcG5Ljya1KzBk6YSS
N+oLrDR/Yokk0c6moMXgFVIYNYv07Uua/zx1S9hHCzXBwM7BMX/PBSF76H5ULU4kFcs0isLsjMVh
kXEqypBhzbsAeXip3WnRKtoeKOPUA8B93ehnAStBoM/zA7hdTjqrEsEpZSwNE4Htk+NUHAk61pcw
7hwycQZFyQGYfsgsF9RbC6GwXYvl9EnqEWKcVh+VW9G4bOpRe/8jMvzvERz9tVH2grOXqUZqw4og
eP+HCzZ2BOxkhFvGX8oF+FRP1e/2gQjC9jqcmbOOCCiWP9nVJe5fTaaK2LVGolINT0+gtQTKB9ks
RTbZJiY7FtrRLqNAI4Y6cKVKYzcPiqi+BuZ77soTjhh983dM78GdysASjlvl+6ri8b0K8GUokPxx
K6w+ZrSNlQDIv0+ID5HPkvN+guBrP3QlDXaQOcFSHhx44RyZlbPTR7ctAJnj3dJ0D5NFlln8F501
Owhpj4TaViQj3CGUrdm9FSJSLS71I6/N6+UyRPvY8quHIew01M43ZDNFiPI87HMCozK9xXzR6fRu
nZsQamR5b4DyMb3rVNaNDl9XcyWnLIvTE1A9AOC7GSiySV2fXhd5hw8xDQJzKi55QguJWH3/tY3e
Aby7EgXh+ZH+e3Vdaj9phi0zJMU0aE7zV0KI9Ar+wL0YM1hW8yr1aSJaCAL8Vcy3OheZa6Gb3vl5
uRLyxOscqKSKOAc+h/Qeiqd+SHNYBPeIeBm08aDdVi0PsbnWjbn7jECsF7QK4Ns7SA45da2+kMH+
9/x0kUFm1KneXNRtCohnWZ8AG6iUmd7Kfnr9ydJ2CLTP//AwmTimiapJtBw5DojFrzkKcjgEuBaU
27ETNy86IH5YMiV7NGKIV+0oe5FAXVRu0HJ26Qkp5DNyivZUtEi2ulvjEOD3/7DgCYCm+AVcsVkN
MqpnqlooY/rKnG7xipX6MY4SEzdvh5BdP/sgMX3eh2P9Gli6+9q57Lll3RMr9S6it7rQJg/B3g6t
usP0gcF5iBTr3o0CaumQYmq7iO6uGDiEZV+4LgNEDG39ITbHtp6983L7ZUaw4NxBjpjIwyV+p5tU
jolAaXV4FnayT5MT4QTLF1IM0DjVLoec8vru2mAq35tytDJFyS2B2hVFIXZVvnAUtYylHzrxaHIP
ZjeICCV51oeLBmXHHmSoKoPLvNXpbhH9MumQWv/8QZtoqJnsTC4rMgPL0w5wb7L3uer2YhRn4Mkg
cOiDztzm+LM0FlPh5367GGz6yb0SJuZoPH0ciYerdCQFKS6SLvK/wG6AMY8VJcfmC5cEh/Zoi1He
i/Pt1xYTpBRv35ItgPKMsB5G76zHMLXnJ0LmtnKEtpOAQHdIb6dbntfIJ5YZdMqL0sHbWhKHkY2g
uDxWNgBk+ZHGlXvmk0SP7TU32orqH/iLRMGRiY6idjZ/P7yAAE05J3Lt8TNy4lKUqV2+czPkc/UD
I5v+pndV22qAdviWGD9AHstJCqfJvR1ppFvUfj43Fv2e/geOL9ncUOrMxWXQpBayJ00qUGMCYxcJ
976he57HLYAFUZxC1nMHJejE9fbi2DMJ0nxBQMFMuk2aGS/2GT8H3EM2aDC3gh8AKBwxD9+Oq/Nt
UwG9Plrp08ovFUUQbj8aFmB3+JrBeeOsGuGPfB1N8zwfzml9yoetYElBHomigDdPjlF/VS41r6Tv
w2e1my7QqCev2dCyRCKaJ4arlR31pJKR3Wx15N+FLm0tL1JcE0MsNpDTG5+w9SN3wUjhkfhKTz7s
lI6I+r8C0n5gyvP8s/fz84pUEoe29znbs2hiBH2J0X3PFYSMON1uV0QZyalnJR34WuFhSa+GDyYM
9oO+EPpYaTsOcpThTlKv9qIS2mB4rIxd7R04rtzb0aHKwoZCRhvR4n2wUE7fsilc8yn7J4Nw9g79
u4zWoZSZd44FT99zNy2OwEmoAxnSutipuQN+xQu9W4g/58yAVXVBOqdRb4X27pu14Yj/ToTLf40C
Ys2rmIx+GrhaxQ4aK6tPOkvIW6OlRuxFWrMPoYja2EtQ5Xg1fn3Wz9kKlX7e1Yo6VeiPDKj49nic
+7Ey1/mZniipzKn2InPELNSIo9BCTavEK+keP8uGRSkEkebCfsZKXjJLESVy4+HPDxfzkOequVHR
1Am+/d+wbzBvAOSDypK7QDlXxjREcNAwK+d14LmflhoQ7XZ0KNElTgWM8WsIS149taKE5n2yvFuM
R1beFPd30oEEPG9ml2uoU3bbEGruGWrJQbbz9uSFBCZyO0G4n7A8zhcg6s8pwEavTiIhILIvCAOl
QxV1FSlSr849l1+RfCwO6SfBW0MVC2kQyHJdXYCJtLy7Aj4TNU0HMzaY+AdYqdS8fxUZ3dgNTlbe
UTpfKqnEFb26lLlSoWpwVv7vJzjovDvyv+q9Z9A/1adtp5pI0rbzVk8FCto9LMujykIQEjPrYf/8
yxWenBsL21Ln9vxzqNy4U7gJwBW+2AtztdFA9HD+qRq4w5+2FeJC9HRi7AtMroV/nLg+rc7LvB+Q
DZ6O7YB1iD6xMNV1xx1WPHHFJxiNfGfD7jZJ8/spOYfIBWxs5dcUFpdrTsZ8rc2gLV32kWT9QLF+
pVm2zVePR2Aty9zI2e3HpoRu5GYdI7wnxCXVkojVoJESuDjf0SQCvbtbnD/lam2hrEbft6TApdUc
5ukY70wD5/0bJmdKBgWSga/3UhTm+vfDR+Y/9qBzx+ErHRZF90+VrG0/3Qx6JsmCUEY/R66q1BLU
itfXebMR3lOG9wohLL9FvRPWkftEMI4bfknOSqtSPi+tPsCGZH0zwAgCwLKXhY3JRLXoJkSMuq3C
TK8z7B2OMieVnuo+MC5w8EbDTcADehlF+BfjyOlbpD69FWnp6qrJjV71Pppq36m16r4pCqxJXrxN
RvwWV1eyVdeWwfy9J06pplCgGEYvn/cq8B2AHB9vPkhf5XkhorjxTASxHUTEAbHK0h24c+ziuRXG
svahhRM43WsfFqByUDdKprhgO2r4viLHNLYzzdG4RuZ+/RSH7KWtG8z3SugRtLX36FuGe++n4bvv
dYETGGFQ0wBrJ1cbr8gYhqhBXn+nEzFvMypesOrlUQx3ewh0XKEByLeJU8nsLnddtn2x9H3JVRbg
QCddPYyDZA9kOzAIX11UINZe1XLbhTjqOeT7FRH+S2r49jmb1DEoeTvhQrg2Vd7JndrVn0V1mmKp
NhGIBL4iJVAmjvGYA/fo+b83NNmx3Y6E9DR+Cj5Z6YgHnDkYQ6UUqM5tPMY7P0Ge0oJyDF2WiELc
g1aMd7pPW7PgKG5x07f+jr4BIIpCT1ViJf79gjN44uU8Oe6TIn/dq9JeIfxfxyOziD2Omzno97Pj
llAyDyr/1vJC8TyCmaY4tQr8sHh7IBJVi44VuZME91u8QGB/CWpLisdgdZVTWIqfc2cFVLRgTv8Z
P3qv+clLBVLY2vHFZFaN2384ca5ab2Z1twr9TZgAi8uhqFPdkBErftUBaIRwdBQVwyIJJwPlW+HA
b6+/VXF14SX0lnAHKc9Ecmw1YRzNOKXnUK92wE4uh1Dz/3ZQrlrJAxnzU9ZBOdPsCXlNZFBs9D/b
artXNM4cb7kLRfUQUGzfKCvxpOxX/iFmdUp6iPzOstbXhwlT8J2d1ht0cNxMaLSWEH/qDqj45mMO
vK7OhpXR7EDwlbCsJx6Xm9iFDN+undKpn8PpmQ9ZsqesQueZBGO7tgiFWHdP+1WaLl839nOHC0Iy
tjGwVAPDAf95MSBb+jDxGczuDUiZfULkxwRySs6edTxbZk09HsJ383k1P2WmpjfYH6+52KEMffrM
AMdv9rGogdazpBA3L1CbkxKepufG1ltuyoVoo13rUkkjPHwe6jgXGsSxuFAs+fWoqcNhhPEW7PyC
ZwnpsQ6WRSKpwskxqPjXpM0+U2PxDRNR2L24StgqnVudSD5oKjuMJMJVIdL23EpzEbCJXhYMU/qY
B7n0UQGBZ/4QZHlwSeLdmJX/YapqWsuftKpmjlULdCY8CSWjFskOVTNTnm8v7T8KYALiIk2UjTPh
zvdrck2kBpj9hOTsIyRypeTe3PGTs6DY7DEDzwvGY6WAd+mOHjBg70FFF+EhhTQweffJFDvhYF3O
UV12xC035XPzekBJTt2pFKlc0+bGyiv+TblWEwnhywbqDeOiLIJW2y4BCAPY56fERjUjgBtN9/1r
S1mPb+zzp/FPGe/bZ/2VCpBmYJkG70IAmHuCuqUB7FJHeJW2BA4pI5pW7W2tS/ViPwqtGP3ioBIW
3F7YGiRKj6IfmC+yaG3GH+ASePaEn5/Obla0D0+OBJRFE81SVrYNospttcLtwMhRmMYbXw3WzQOM
sQKvkvGRmJtlXz57prHrc9yHz34K5+M3mGMpR/XRW9DfsthBT2DyWFUywHChgQeFxL081W6HbrIp
O4q1uv3Hgk5RL88q0KBBnghLT31Tz822unWXNdAtD0+z+AMBkgOA370winRzHPuLHjCMnLZZ2u6M
9Zc0a9TreTm6BsdpLDJvadyXQ0/pbuLV+NIQWwXijOx3ESnzpl6W9DM2Z9pgCEcrdYANjdFAWuu/
8oZeeYMpZ/JDWQ3h7JPJkTO1NKZstaEIKX1U3GtfiAlipQoYM8+hhad8Oer8qK0i4lQii7P0/wXx
fOHCkow6/2dhs3jMST5n+MVbewD56K1CKn/z7ar0tZNTPJVbfJaidYiSj3E0b3yvjZ0+PvUrKedS
IuiHZcNyj//Vr6mfMK3B6gx2wQP0x4N8YKYvK5VbKAVF7G0XvNdB28NNaXyTrjDhaSdZabiKDjBT
Z3+nEgl9TjL02mVcpyubym91POAgWnB6ca8q6Jdt1Y8KOoJNTq6wJS9rq5Pv+WHjeL8mc07P6Rpq
eC3fqacOcjnDz8/nGnFvxkehqFmOAiUDmVWnp/0liEw+2KqE042p7r1Kv8Sxff4xtRcPbU8COslf
hJSnZzyXGQ/WaEJMPA1meFOLGIr+iaiHHbYlnlC86XODjsnhr4AChc1rrmpqbSHGtb5utNbxEMgz
zBHQZ3kwfhzYmDsLZ7CBcKH28emDc9kGMoMs5B7RHV29IBwwocgO6fF+HGeZ2tvDlelbzYZls+DZ
1DDvOitjZXiJFDI0rVzvl/1ZwKL3MHRaDiljOgRSk2sJp8e57tuD1zeHhLG8wer+UzhBYDqq7qcJ
MEenIvjrctRtf641zeSpfSryuJ25sb8HcaCikkzlraWH51VJpeWmkTZzHVKz06RRoKhISEGLVYQt
4VnC0XD38LkxuXRYOKRwHfLnVMawUYNEoLfUcGChK9Ab6sMuqdqjzos4evL3B9NyNggi5cudVApd
XG77u3WENELNo5ymCweTv4n1wxj+cxxrxzBsdLp1SewwTyDePQMNmi3lW7mt3wGiQc5faQM0Nfnq
4REAefplFGTv8r5El2fOtMoaPsSMY3rF4XmT2VBrpwdLOwIu9Gi5BPCf5bkmFeN1tzYhW1CBTATq
E9Evr6M5sjLmD4bNB8NjUs56BigEsVuOBWUOv0sCH/rD5FZ9IsqKgwpp+l0LaggCH5EZanD4ti0Q
ySkyi7cfOrLbCFOKvkLnCqkhoZ1dybsPE3Ooj8tDQ4AIQXuOSz9YvIufUeKhM7NJJNb0Fnl58z/C
wDP9aEkocYyCTlY7huRP+/DIkCZ/RyJq8aLPyri1D0zB6BgIi4lLiKwh7qXWzxFpfE8/8BfiYvwx
pKXf3YM3p3WYfbkZLdAFnnD/wVYalgAJ/Y4PtPd9uJjpvMww2d4gHa8goL8AGsvQ3FBVQKdzzF9G
dIJ/5MG4+dzd9Oz0Ke3tD3Y6NlWYCXjBl066QZ///TdCYyqPU/UHqKQT3exrx3SDr6sXv6Cv/9qG
entPFg2p1NvlBqAHpGRUPBYLS3xFyyB6W8SQm/SWyhOPY3TQY4+jq4UoB6gKriJlaCmpVMK4D8t/
5xjo1BQNGpnINApkecffRabPQfWrf6LlKEupUaJ8dGKKP0flsPjt71PLUxLfuz4rL/Yv4EcOFEmX
XKV63FuqoaK453rmSqioaMSo5BQ/1T+K1bGH9P0JMge/JAk+JSgJnJGvmILixLn7YefKPPHCkqRb
fDDnOHs2ruKXB+UhfP9UE6S3Zg2MsuSqOyFuCnewu4OIORtMX2fyzAdgobEhNClmiKjYH32dVJqm
TMVp42pzO73hY2aJEU0H0cW7y/+m+JgkgYLwxqoJeFy82XSyNRg+W+8Lvc5h3HpKKLqXDwog91Re
ipjrRgbxE3YtZPBPRWgq8xPxqUOFd1XvmHxtojEBtHFwSsrEJQMdoaY6JhCWDCLm9qgeLCnmxnij
CBOEnkeT7Kvj5ZLPFWMO68YkhxHspLC6wqVY0e2DNJkSGX8iCrgFF4N+atNvTgyM1OsFAKv9qPbV
vhUhRjbwkjAxnLILQ0W66UeIZn2VLGHSJYnkpij4f8iUy1QNIXFv9zjSacyU0p4L/aKOkvoysEcR
FmJssQea8wXawy0qNHgHwlhL6JnF9BWuCG9dKO/r4z78W+GxUpEABM1oAZ67r/gnFytwkdIdot/C
3XhnB5rtCMpiVBwG2oWrLGTWQ4jx8fZTF+KwGZ9z01uQn9ZoTkd+8Z42AIyttXAXapRXgErMp6Cq
9nteANbuevKHvmuZn50CAUZDDd1HDe+No3UHhrO/f91UD+DTuI+SZ2DaZLqM5t6Lqa/6CQou7X+7
oFNHhLTfHWuyVzgqlRpOrVJ/Jrhewp7lR5kI9KXmaMn4fJdp4Kmu7q9vir/xodfKr3nGLaYxUOkH
nrVYr93CNI/PfVvG7y9YFWfznnpRko6oOnS+bFYcKLz/0o1NL5uOEXh85DbUk1sQ0tWLijnt2+6S
3R+Rn5m4aYosiPt3z0i4bppgh9GIUbjKOnpLB+us26Ky3hxScv33z2cFzkJ95BtYZOstZk6rQcaq
/USF/JgGNHYAQp0YiV357UbQ5a1cR0HSt7XzypAK8HY97QZJnEZV2PSILoMmpSGD0ZhVsaMaNITI
X2joVQvCBK1C2ZWPRh1UROnWy99hv0sg7xwnum82jxenCUczs5oQbXnMxJUIP4NRozSf9zYwp0R8
5K4UmBM/pmtKMzCZ/YhH1/IXt6UV8gGNMdYmWOMDpHDi4AuGFWxwUKC8talDG7xaa0zBgbx34QLq
LJK6f6l6/+ThQpcmqGgD1JQSNL9A9yQV09tw94rpoBMuIb0TZp2jOmL7ciM4uh3RKBoBXBDJ+eiv
OgrmcrEmgDYYDQSmXlyOuV8CDYz3vJiwKCJPRHiUuxgIjbzvbjeANtcf4PXXMBPqhnZfL6HqLAis
M64jiLlyckFoH5SecX9DHkCnjQwgVx2OXoYLWWbKIDRIQzhQ2thRHLXPRaYyJMEo1eiqJowuq8F+
OhJq+mupmIF6kPirb/5lMXM+VRg3N5Jlsu5qbSro4RbXkqLUhbpzQSe1Sk7Gas6/cXQbkPNto1+R
N8M4xoG8/MuL6CoPYYYJ+O8VI/i7D66+HuBSI/zhj4MjHSnCiP3MS0aTYHQGhyHbivwLdkUoanNX
hQJBNWEwQbM4BJ/FRLkU2gQOuNYeVll8YFn/gFT99Yw+F9LYZ44/8ixRKie2R0n85hwdTAUqbC6C
unV6hY+RQFPBsnQ7/EkM7bUOuB8dNmflbfQ+IB8XNkD68I8GTm5opLZKWSA+VOo2ncpqMoFW0CGG
9b4QDAMMXbRWOQj6bjw1TatC9SseCkGRdttEXIHqtQq4wQpwkCa8nxYP87g5RTzqInTtoUo2FXka
4TOQBe8Td/i86AHpsd9q+s4HUb+td7PQExKnTx68VDL+fbgXHocPPiYcs/wugZOUB56ZuNvR6mRr
Z1+aZ/IydTkS19UVLB9Yi0XvW5pd2+o/SG8jtrZ20xL1NVi2BfkjClRwx5vmapijCjd8afj+4MMb
yNdRG0AIzoqGSxwubRrwrQ5D8aX6qo/td2HOwMbEzG09IJU6hmMzCoYzepr+qExuWd/Lsbl6oZrT
+1TKmwMm4V2F8GRQ8cE3gIwAfUC7eCSD327/m0ooyLL8HndMC83uUkAk0kPFhGpaUoDpkkuLw2lN
xVR7HR+lOXEKo0DdjiloAmk7qqx3qCXDEGe+uzrq41r76UFYMulphCMpVEhL6c5dBLIncGHSyzQ/
L0riFfzfxtspvNBVW8ZIjDeCf8neJMkaL5YcNZMc0gprXjnSgFVWZnBcQoRUPRVPV4CVER20gcQ3
Ru2ZqRPUkCnaDDIzud3+nx/YhyesbANUYpNxUsg3kA8dQxUPW5K8bnIkmDxTEBLKbNF4OsOkkGGf
vg6trgYiJPlCJv4KVyaQKi7FLsh+zITnsD6gqvORRRvXKdRRXgi7zZbFUJpZjeItrLAlzTtoltGY
QrrqbO/hHgxdjI89+fmaAz+a8TLb3Wo06vfVBnpO3Ev+k7UgK9WU4Dfkp/aF0twzh0N2OY42F/rf
MuK2dWLdEw9tGwx/CshmQhCrAbLey2vZBN85sWkf5YJdj+Haf5a8ba74tOM5rfhNSyPT2VMX3WID
a2NGGwNHBYIyGQzAZTdc6BWwszITT5H8D+J7bW6i22zbL+5YKaytmWq6d0RxHbDAUxGKo7Zexbdy
Xwxq6Ik50aj868Xs4lOI+MDSYCTUYMbnu0u0mFSRGf0VPPnuZ7KZafLMg4BLj8Dphg/k77Tam5eZ
WS51x45ReVOEf9KK0n10hWIOHHym9S1t2sUaFOEr8CnXJog9Ic6bMARuxNUtV3uhb39tfNU6kFMj
QYQ42yZhTpcd98b+C/O3xrXhOBC7h5HJdqYfPZQrPDia3Wn18At3GQOsjuZZ4StX5Ns+g5ciiXKe
CHHWEZrCWU966LH8IrI6RTlgySShsGBaG3ieKlYjbjFUKse4nbmvx/SU/whfcckSi/tHMFr7iBRX
4590a+Zck3XcccRKtW8JG9Qa5dl8dn1p+hEk/2Od4ttMToMlBvzfXB3rsBCAh2F2s7R6D8f2Xeky
Zx5YO5NgUtcaczF4IAEnDFSZK2A2gRqjxXq8INozEUqi2sUUquvj6jdzJKdaPN+vjKLrAbeO1rM8
e/Ch6vDD5A0Jkwqnd1h/wQRdNApXcPDEBfvBPblSYEPU6hJl5cZDoWhbXUl/OZ2vl+uR8td/fB/M
Fk1Nvd82W9BNKhOzn3iSRO3+p40Gj8gEsQOoLarSxj9nrr/8W1Ka7Ik39VHkU/rz7BGVHYaNFMwP
PHk60GS1UZdl/cMljVQ8y3DcFVFpQD9Ko+Mpn/TnRvq1/XmD9Y5AC20LwGnJ8GSbeXulZZ3w+Mw5
q+RfhnZeuRgdBzILRh2zZIAPfZ3CqK0lvFW92lHsok0fMkecvFJQ93kuT6Ngtr0u31a1LnyZlx/e
QgAFgVoZ3BBIh9kvR+zqVpB0rva/SacgqStyfk/k9j/PMR/W53amWP4dAm6XUWNOZwCVzZs8L9id
P5dZyCDTv8GKqjAqJ183J4OJYi0FhN9Ev4sJEbnCBwQswZM8dcX/hAOkgByesB1heoP3xp427SF2
zsjXPG+E8lTYMnCDusbYGWvAJRZBaPCstKK9FdyAtyzup8tu4VdtFcCPq399cIDSM4vjAdoULLa9
Jd6pAgTm3lNpDgH2+TxVVu8my+1Oy9+O0PsdVnEQrio+JwdQqaEpR24t+PdEljou+1jen4aB1T9B
Wm9ezzpuetCudxRiV+XR6pCZmiKxtp1ZX/4I95em27nK0o2rdassV/MNRNsWDEHy5XXMnA5mb8Ru
f+ns2dXIdfmoAc1+TTde3APxp5Ok/KAhXGEuJS/w9yawvIJnMyDhUOr114dVzUEmdQH7xHu/tUr1
VeeoM6Z1N6y81b2qswpKTO7R+dw6LI2jIol25NxLmAdUlPYKFQ09wYl0SBmscCWNZCrQm69OhZUO
ZWlk7TlBeN0w2urRo2Wu9Ay60VhyzErXFzQIFo4DTLflZVXreQDI+5DpV5tD8GaOHEay8hU5OzPa
fGaeSuxNirV/ZRwtgITWmMQkI+O8FMj5HWqaQWX3L4x9N6KuWWgBxpW0oNqS/qwgZ7MJmgswv9YP
ljo+rM5zCkz8xnhCILoQTNALwFZnYQctDkvzxgkvhja3LvVbqqY/oGMmnwf6khD4xV6cDJP96J51
zPYvUwDXAfhJH3y+xHyYKk/mOGgIy3qOVOLJgO3UF9aBvbx84G8jKBdy/Ro5+cF8ICIaPg6rIJRG
WDlMrcc4J6WESgjT/Hzb5TtATYMdZvoRduXXP/VlnfwevN1ESULulSId5gJaK97N1Ky5yaHZgmUn
zrtQ0BaaJaGK8ZzMU4ofDSlzWJoBWDCx5dFx/nsDx1KoBd27Vs2/tf4PeLHbzhIl9qgG+nGhobSH
4bG8rXFSsXVmBKPCEA3rWH2qE7uyY76vY2f5Q7+XQ8hAfiNI3BmC8+q41vkF/pBqY41fghCVSRdN
OosT/HRAWr3/+LENH6MFx5zs7e+GGMc9gpkhal0UC0pJ3cqVq6fGzvXzTiH+RR2MDH/TLrS81maP
EQSb+y7M0sI4wodmnroNcFyayl4roj2F3KUrc/nT8PouMbByan/ytvNNrfDgIogdI3Ndr5mabff0
hgeqIUAMxRhO2y+vu/qXfuCL1/ZSUWpeeNqxNp+jFsA2sZbStDJ75h6aBtisiR6qWOmHvfeFA5/8
9uD4fS2lAU7/ptO46kRaE1LQgtaNie2bAm6EclCLYDnt0OKpN4l9Hjzae48FUw05jjslIZFuy7FG
wxxyU0R/pQPoUtLQZtoqTOd1Hy125QFsZEfCpsgE8lcypAuuqtzSTN/x1yDI5gEIbyI/yzAzLYXk
GCFBIes2CSx4Fhj9dVpq0GHpDus98CAS9OD2DVo7ieGMKTa6QO89jqKqsdzahyoShvwR3f/9ZswK
EjF7deEic7YBP1guIWDsOmnz7RL/WURhmpVGKf5wXzit7/lGFCZpoarSu4EWj9ne1u0xHfMkVV3N
2oRnp4RtLrTiCG2HiRGThBnlZldrrHOPtwqTHjPWDupXQZwq8OpctVWHYdL3ZZ2EgJ7DBnszTbNq
RSSmza66ABe8K+qKPL2+QzPMjXup0eJZmJpYrVHjCJQfanjbq1TGHCVOIiirqSmTMEm95SdVpgQT
EcPvLmSEvJvqjejGJQwVMnIIzoIRx+azKXWUu3ILIIgSWnOUwtW91/IIgA5aijkw4rVbKV5dhlkF
NWCOd2wv4K9WjlnPbgKhGRix8J2SnNso5S86WLz86HdKAXWF6nPQGT0IChYbx4ilrt2LD0Owi9ik
YfNM+u0OAiQiecXn3KKatqtBAPG9Xls7RcWEeHTwdjGFSMezlGBtgl7sdqyuVtbnDWyGiwCKlHWW
mH85Gh7WUwD1jExBAUoG0WMIbOHosLf/17FgSEV9jHkxDNHVVRu1+6hko2Q3aE4a17X9XiUP+vIi
vo+Fzgkf1K67SPnZLLXQSP/iF402IL71dDN6xk9IOVB8ELyjjZRvjbMwI6R3TDSGceIsC+IVTuA+
jDCfjX1NwBOYFru4dMWiFg0YJZ5ZSHJFuo9VQmrmB/6nXJi1+R87B/x1pfLup6OD86YQtlIHAYfo
6/F/QMuOy6p7wBFzmSm0vA1+de7HuW0iPFiZuBpjbCVoi2Y+rExA1JjsQrwdQhk8hZj7siN33/UM
Odc3ghUBshq9mNgJRVkOOhORoOD/gruJBfpLSdsXCnR6GijGnY+KOIlPK9c2uH8FXPzCKNFmvMH1
SfPiof6HtsRF7t7Tb9Lh9EG+nI0Z41BtokcdjvF24dOUdhRC+1pf0IEAT/UrG4Fp6CceAzDHq83l
mfbAPX9Aqcs8sIrhVooOjpF0jM5zrsxyTcz0OC7qtojo9qvL/hTaIrQxBgPemVNGUMPslueo3j1I
onKpCBGKrQ0E26PQttofYrKlVl4y1UXHfVsQLfKeQ1/Ljbhu4UjHS79LbEkrjn/1TYgKvwfRgyr+
LfKKfYgvvtNvyJkuUGpzlctSZOkadHbBKK/rQxKweuxjN0cWETM1HUJkmRvFVsWZbcIshzlcIsIE
y6KDiJgm3w7OyOVdDBdrSasPyAkMW5uUuNeu0w4wbq868PBig/qqbPUyc6XN2Ms91ng6d6zQFmrx
OkhOfZUBlBCaOOdocP/JeMplpQ2zdnhOtf5E1Y0+R71K/P6tSKpHOSDVdd2EnqraDa0lG4/z7gUS
u5CAvfjmqzvYRD7BvMYMoK6s8wZNwDB2g2cZ/JqO+y6svrGzzbyB6RRmytxGkHvEHw3DMspmonyI
i+ujsrSOhC4TrKfpp3Hbopk5qSc04aIwIsVgnMZvgGlLlgaM//seqzOO3nPj9+uhCcMZG7/XJxOQ
0FPp7FfzdtLWba0OfdS41k9VE6F+C1aFct5A2bJEY1egJ4mGW0eTmKaun772h2LA/JJwPXGT0DR1
y4d88wd4dE5kd46sWdAvu5wLMkRG17wEeLCsdr8kQj8jENw5FqBz72T+zo19Lt0evQa7Cd36eQjX
AbHHQVuBXvaJfhVI5er33clbEKsLgI1+vijmkNqHc6aLLPHsagJvd6CrKRa22/f4xSGGNcSnKmD1
rMHg4XsqbLKLAOxx0byN6/uGU719+ibvyGTWTmVtrUvPN2VzcRJSNpO7d3ey9c9s6PVw5jRVsDGs
TJVJgm0tMXt06NzRIhLr7iuHLHF8ZlCWGKgf9fFvfT1RlfKKhsALCn0YUjUKWvZFJPQfrltf1ZRq
zVFi6Bd/emoivNjQt/Fc2fivOc9ZYp17s3Dy3EofF0kZuQ3vN+QSdHIRIQfO1lcP5P0lBg2LX6uP
furx/s3LDoxX3fvINRp3L4VclineepImJ/QPH18VhyHRdWji1Jus0ozeCN3w09x36C3lGPX5NwVE
gBC836H9LYoXtruF94+wJzWwXX7sYQlkX85PAhBQWRQgJhDw93Kh2pq0Yk11pjEZSdchiPyuskXC
mUzbVaj16StEoc2ZerA1NPKpHn393m/zdrdtGgIJBM2iIyPzpeXLR8S1NTEkRLmBXuzP2H58iv0e
cy4wOBvDFAGHIjayY1zOwi1nqnoSdbd5Y6YUE4xMBGfoYVAFBHv4f2z55XNxnfXdemA747UN/2J9
TL2hwVQr1RjtVHyphaLwc/yOgLuy+RLVXqMBAcfrPt6fhmjH6LkjE6l72sI6sDAmku5axbJrqk/5
rjQdYlh0883SzZeX55DFsJHJtq8AdoustyhrMkyPhxsFpxrpSOHnri2FhvuJwSvixiKNCVP124fK
XkgtnZoTqX98I8HtOgbh6U75TbyoYXCJ8i462guiu//nVfBXzRcY9IYRKmoxggayD1rtWYi6IeN2
o5vravDX9qvPHsKuURb986auoXNxm2C0Ey9nRtNXVktXjryZ292L57H2FOhKc2DHrFbjZxku/iom
W0xeIKnwDCH+V2n7m8NK69m8oJMflbBtT0EMIOY9EK5JGWlUMPcZJcZQPxa5H1liPTX+S6GcaWOQ
ZCd+k34v3HQumc1bVedPcWd/m5KP+dXtGjUO0AIp8FYCiSf9MGWeNaHdAH1zwWUQ9cV5GDQABKlw
XbC+VKDUyIW286gvW4grp3cz0NBsD3py25xVQM3aFhoQkFGI4EXWko5SVLN9u2GTPG2ZL6X7CEP7
CyuyNq9Dtt7nCEiqIEQEgS6UPzCcfoHFyQd428cy1QxoQEPLkGH/U9c3QvYySIL1OviS6dG1OYFU
ZC1RwAsHOkAhm7iwWdF3+b1Wi5xNFhI6kxcVHwMt8c276tKPWw7TvD8hJ5S5oAtSsD5Q7kKB4135
2d9jqp8C2ph4eO+8xTt+XbnEbob939VWsZbAIIqACO8q2qn8NtHMRYgBozNCAmf2g08xAFIrvGev
n1haV62ASVJPQINZ2/5SP3R0N1zDHgw7C3eDhkBivhAzmqYbfwT5l6dY9KXqJVcX8U7HSlGU4VuD
/q8EC67/uwcqFWw07nUqhiNe62i8gJct+wVrLb42lHOpmmSEp/Si1vTOezlumECSWpUeC21Xs4Wn
ejxglnRgCpZIKdYFn31WFERpRfhfS+3w+7+oV4X3aWLUH4+/KHbGKaRRBSq2gLQtEYJIux/vW2l/
l7BFJk0FLlxzNKFxmvkDA5C98KJThbrbbeZ2weSkxMsn4XsIQU4PtpATiiA9OZ6FdjgdU/EzxFuN
N+OrlnCfoUj/ZCi6AoAwrCdFuctlu6XJvKJGfYyadL5T+v6/9UAvdK8c/1I9sX9iUbqwP4boksPl
dFDtQbOQGLYdO3cAUJ15/9E5vsxlZu3GnYfr3Js+EkplgI7gCad4sfjCfSPSaNWxi5P26L9djX9Y
96FGB9Ux8cLZfAAfxJmE2nxyRNK8Tp7cPUaQKDtaJud1jNZwckSjyMzp8T4imgaGONpj4XzLf4XT
LYQMPhs6FZ7mnQcWhgdImLMwDzpyXJ76DpfWMD0vrJevhMCAOzxyTJe63jcgZt/6FFUQhJLi292u
RDqRs42QUGDXvmWwCLAuLQP6uGeVIGexd91Dz0BEGoVHYmmbnicnrqZNPHnxzLJkEPSXUCrSWoO3
o++eXY9FU4z0P0hK5vqa3azLdjc3zvMqXiTgf7ySXbw2+7doxKdEOcVWmiOx1/ypeaezYWWYoGAt
IyHiI4Ok1lvnxRbX04oykXlajjf0g6PLElzFlzf9pnO7JDBWv4m2EcT0Qoti5TQw0egOAkT5dnVW
XEElUI79eB1hF5MjtrE7w2HHx1cZC+3S9d+PCXP/O8le9a8wiPc8z/zX3VduSgStBk+P0qEJ6FmN
eFyY2bujnwXbyD+gJQ+GwlizAQ2kCZIQZo7gq0yRCEGG8iWWmjB58IFHZQv7hpPnpBlHkCAVwQxj
kSwAQ8oRKfRuSv07XCgdykWcW/Ios154ZVnJSAsXS0b3/KPGmwt2Z6t5Qu8E2jTsSz28WthATpQH
WISb12GFIOqzfjIkgmYiisHeCMuSUy89TfE8aRSagKwpMXvd6wTbwMcfcJjFaTuiF1DsCSTjzcNl
C298DQY9bTUgQ4j9yaXNccTmThvE7PDyGuvjtMZ9w6c9HdkZnsGH+DUFOjCNZeK9nwzgUe4EtGer
qIGyOWacINqRj9Na9zfsmM+pqlVc272P1nU9ZnRTfyS2SOr3IoZJr6oDFNrV6AMuLhqlMXck92GW
GnSg1SvMT6yHck+r3DJ9tOGGWVBUSV7lIxcilGdJLT+sSD95HFgPyguQMT8oXnkIXYNwVzFB+MWw
DIP7MkpGf1vliceO2xw6Z6upsvi0ZEqk2NJOGpcxDab3pngrbQZHwuhaY0cET5FkGRckUZd21D0P
RkYLKlDE6ybumxDSxTyaZA7nAayPKNONGLvFSoVohLzmsrMFqERHgVHbp+HgwP6shWBuKdhra5WO
k+em374b1jvW3p3ccoaYS8SjA4YyA7VxbtyMe2u7w5ch13ikELXPK5X9j7emRN2/6dUC0Ro2jBBg
2AE/TULjZp9wEzrxevecP6xoiZjYc52tMuxqEP4/vi9IlpJXlNa5gLSWR0cPzPJr8xmXjTaiK5fr
zpYs+3+0jqyomln8doAyqpvwy92SvTK4l6kXy+J9bnUkW1q4n0AD97lj9fwNwGaPul96x+yGglor
RX8RTfzDTmBGb2w5CsZOvOUCLGSRuAy5uznxDqlKUm9kp0hSTv+QD814S+5sX6qSbXRtx/Iqmhrx
mQZ8ushzPlYSmO1T8gKXw6ZVRIMiGDXPmTkzethAeF89vE0LGMnpU6ly0kvbPRlC/6cGlkl2ZXtV
YvzLQjgInQqygDsDTL02B/45dKRUWZf/sdygFXk2OS7BxlgdcUsgUfyW+TP7mjjGaXIjZlFgktS4
kDJ6Q14//sdObbDR1+3qVLY9QyCjqY6DUbw8hO+3w0p+PNU30opVGsZkbp0ZqGR/XQc9oVtn7N8r
+yneT4EYLpKoZwyKbYYi/X4SZrbqNi+fAPs9hyQRldCCq6Rib+EqsnqUPJxr6gl7VcrAbtrE7dQk
x3tyYkSXXJ2m6QsT8iOqjsxtcuezfXKO7ZauF2TGsaOVXzlsO17ce+aub2xxF7UOalebIZldMFVU
HtbdTdT86mlxe/P73Yjiij+DVdE+fyw6qP1C+rzMmVrNV8+cQdqdX+oFCTlXpUUsJchWaOMQZ5xJ
xshz1aAm2g/WhQChj4Tu8iZmtIK9pPVxugXCXgxhDRPgUtlaupyegGNaKIc6+yGhyrwJlh+HgcWI
jQM9d3XsFlQmBvQrciVNCtGl/9zeU+65w4a0hzS9+RtpPbOb50HB2KJrr3whrQhidtRvSJYUSxVq
M6SLiElX5H2TyvFb5QTyvdU78zutIgrA8C9//koQSGdKc9zz6OgUmKJ8mFEjT9RRp8I2IwFH0lcg
P43enUksE1WbJKirnITNtbGs1BLryO2puqPEp2SbdXKjnx+p8Iy8ufCyqVMD0j9HghV5DktvT7LT
CTAJpefiUTpyFQCt1jnTahIrOWUhNI5tCyc6B1Itj2g0XemKGvTBqGiOLa0auKfXWQhrw9uDdc3Z
qe6I3lzXEXgFoARzD+UPrNSJVqx9A4JzHeVtU8vEFWYGAiNzGpkFynmCK2QNnvJxz/hp5UAsHqHW
W0ks+imgED0teppaaKyzhN4AJrLfQYFsAtKM4vV0cLDB7Yz1NcgnKU0aINlaDv4/BNYGVNioir2v
EM+q2JpBAVHavimLDGZsXgC7zBIoBWj54Kuv+dk0KZz6rBNyGP724jFHYVuDSaEN241PYFz1nF/s
v9/AoJ6bIQBWKMEDXnBTo5AOX/DvgNh9dm3rZMRjPylvnQ+UiluHN9/aJ5IdX0jTHRflXtOj/B0s
XLe6ttkEYUY23CpXj0y2ZSnKiMPZ5BBdI5wjLhsQMlNEmzuUDkwMGNjMQ848MubiIx/yMdJt3svG
qBicyw9yJBsTVHPh3Az4Y/+Dep13BM0QsO4CJ3N2yeFDY7b85Q6A2/prEQMbte09g6oGma0tdVMH
gFvrTtLi8fAYE8/GazbkcUIc73MW6ieVyJcCx9GhXw7BYi41ec4WRTDzG4V9xujKBcBXxeT00Hbv
O8EJkQ6VLU+MMCHuCwIodaTKC5TofBiaP/cL8cZfrgLcXCbJI7atAZ+WeUcCLk3QepFp+L7CISqg
e8cNhmQ88asCRRLyvzAJo7AdRFrVcovu+FFQH80Xky1uoJho/TC5B2UPX4vTOKqW2lwB3j60+8P8
BBK1yAli3OyMOtoTt/wqJ7taqNBBRs4153BOgBy5HFm2+uxASxoAGDm44XKQtijw1/4G3OpOyDcU
iCMdcMB/5luyATInTq//CBV+OxpKgftgiRvd4CckA75LF8VhbZWzH1Cm6SYM08+9wAlyd5NeGbcD
raSIF56FQJGgzq6Q8D1PHt/GsGHq3S/UI31Jfo4finusOkffB6hxyRg6cTF3d3PWdpHf7a9irqtQ
an1Chq7wNmcUU5jB5lwS99Ti61ZX1grDzxBYX2Bdg7EmvVTy2qAumJo7ZVnR52Go+yQ4+SyxMyTr
bPzaxkIdM3Yq5zXTdabDri4LKCVj0Oe6a8RVbBGP/tyYiOsgd7WWkkyjtmtz3f+AhFxoHWI1fmFT
fZ4Szl0zoj/YdHNNH26AlPUQV2HGG87h+pjQ3pP/+FiVhjOBGJpjMD7l4BTNiPAPI9OqCVqNsyz4
exGSzdDlqLoa7/HQP09jichjUVKQFbbbnlDlpoOmoi/OSDy/VqWudzG1dbIp9hgVrkC8h0eTE21d
SQGjbGQWkHESIymy96rjeRCVzidegcmhlTSEYD3+CQDjyNkjOl3/ukzOKUR2F61CnH5z0r2T3PIb
LkvWTkFZ6xlE4oi6f9lMoYPlaUu/qE6tiWdAxEN04YWTmGjVKRzau1Vp6LgbnETGrWp+iMmxekM2
VOpNcNpq5bZEbNPwcrBBgP3fmR+CECF/soqWEF97+SSkTJ4fQeuUWyjG/ZYwX4TYRkpRwyNERJRC
ltMkmQzSQYu582Ie4Ug90/9bOztT2rp7jM3yMQKc3HfcKChfe740nE0gKWaYTg6LJLYXWEHqPs6L
Qw/yFzrNxQBX1apM43xgrH2ryYC2xiNYbExiLh55JuNDIyzWFOPgStkH3QyMY5VHvY4/0SfyVdA+
RX+DWsx2CW1MMD3MKJyoq3URnq0MOaMnxXHzPFGuJo35EyB5yuJGqFTirrpR+THgiSilwFPFyFRx
Fc9hLd/c6KheAUOHrfnQf1XdStF5YOu1Plx0C3bMfjGb8z86j2UZ/UwFuxm6YnCGsv/jV18lSZl6
CADSrfCklfQEYKLtyNGsX63sgVU4LmrwC7cr/Ne4qR7tWeugkptXbfJdV8fIB5z9/HKQ5EtZdcQ8
i4qYbgkRAHoirv8aDHVUIu9G8agi7rMtVnipPLGRL1KUm9Ig095lX/ttNv3n1WPajZhpbLhsYiS9
ZfEDhb6R2q8SXB6zeU/6CuAFglwYjG4rZlQ2g5YOFM09azMJs7u/90Wdqg4cZEN9c3HFu2GLxKiw
Lp+J2nF27OKJJWqac5OBF63ZB7DYEEDlgl5uBRGXo06CUOHIfGftVADtjYx+XET5ufTLX2mZAwPs
GYudHw6Slbc1NSVs1v9ux4Ais718RDNNywafXY98c2JJcT/Mnks9Tr+L0A6w+VQ1OSHxYNQVUBLm
Wi8cLXebKSn11S9vd8mBQMblyuKhLAOsEIv+9OnRDv235Eo2nh0wxEFM/76qA+UGtmR8jF7GnvKb
LSnPsMEThky/hUENlNdEbZi70fMoHEfliwc+pRQGCV1luB8NBIXdS21AWU0wCMmVqGGnpbQoqlyf
X/2oC9LRtCAj/n3jnxe7A7ys1he2wSp27pzoue/e7sgEkUwj+6wC7iW0kwSX+GmiOdNBPJTCCylR
ZfNKliH+8N90IHWt4IEVIlSsx/wxXnpa10SJfFjAmQ3bBsBbL4oCowUfo5E1FfXTwMZLGP2e/UUE
irDA0qKaoqHGLumk79lJPrrgmNLbibYN5Hyi0feQcc9SKkqtf+3hZzxCZLOKoX2lV5H51vyYZknH
jQtvmB5R9eDaWatuqqxhd61ZPi8gqPEewSnrm85J4SgQAHhVsqIz0NQQTZ8D1IWkv3nc5YM+kIGL
B/akQNEYqX6NmujaYMsaLKadjmXBdW/dmTD4zwL1f0kJipKaDc/HxD2Pj+TsasSwKEZ1NaSho+vI
tUgnfqv3BvUmCJa0ZbHuWKFnAXL8V+f1AMEqNWGRmeRO+WPmP7X2XwJ8D5BomS1SCz1PCNSqtmUi
fGtK9Yzm2sXWmW4NVTE1WgK81HeZg07u4NlQufUICMIKlPeSYZ1rsVdVjhI3MLd28TNTFXkg9SJe
mjlrtoYA/xNmlAa9i1VnGoWefJA8qPAJkG5oEN6rpwhXPWST/7nBEVDOqeniSNjiJNC/vz3VgKLC
zniLh5fngz56hVe16ERfwaQqxCtReaXdCcwEFIkIeVGvxQOzJu+noQb9Le4kcRq+pNIM9f/+LsRG
xjOsFvPnK7IhzChYsmtes/tz2askfoFgTJiVSizhoooUvlvZlBuqQsRqKcjziaWNXR2KP96FuG/0
YeDSUqAmRHaQGmzR6rxQE/oijk09VpzCddrQQ9jiOWP30b2vtDhsS0p+T9mdy3OpCNUJa/lsso88
4mD321S91GhLY+6q0uwQIS7XYC0uzAOnGTsnnghmK1n/qVMZ3XwXKOmYSQwmUOSRCBVqREMrB5L1
yXa3tdm609Q4skPdWw0NNAUNg3Pi2VIlp0YZKvUleNfUhHua/QmiKIGLeT5eXKNOaLrS8XU5XaR+
kykBJHhuanSyCfZ8qu3OBO8ishOmP4+wHJd51fLuUE3MXiXmq53JQlAImDbdQfHLtfu1uJW3Cmoq
nhTDijVZ5M4eqiHat1GncCObXLwkXQhb1L+yK7oOQ3rueFFlW8xGKdtQ2kEDiCcvkW3bcboB6WGZ
N5ExNCb7FK/xgQAaKE5LCAVsCbJu5fAMBRS2iBuqRAQ8PGaD6Hjke/KRCs1GVSrCe5uzoYoPvvNB
1nlRXQgyJciCsTwuzQNnjGcDJRNt9SnX+YyrM0CYhi7oe+p/9cXCBgwFPhlKes2NwxRaRtjZnW0B
/jF/x5oam3Bay9oZnKib3ELYRCrpHoQFltUI2NUhcioOAC+wzta4eEskUNC4sIMWRHfnyaOy2Gb5
JsaCuo5T8+aTVlwk8EKeLKG5vi6OoebDDpUPr9tISZLbNHtTnv3h6eH6brMA8KA6ZX3epioKmrbR
qRzOgcek9yzAB3g7Iwq60sIXXYSu/B1XhrjI6UC5KcyHOIdizs0I2z3dP+q/wOOn+uU9/L1IypWE
fm2WCSxr0OE4QZx/ybPiMr6gbVf7DLcJyLEnzTskiyzthrOzLBLjvwgYmmHdznwmikqKLr4CXgUW
wDtWLaAP5/mxiAOgLMkJKo0C0XqYnVlSxXfvlIZ2+WOSVKCP9txgwbhSOR1a83+dEg==
`protect end_protected
