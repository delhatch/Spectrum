��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k��ib#�Y��&UA��?��?�%|A��͟ĩ�x�Yrl��睇�Z�Ǎ/�|���ҥ��6��*�h����l�(]wGdZ���z��3.��)�"Pz6�T�
�	Q�%�b�w��0-`��Pv��I̟)^��a<mOUkyGL���s��Uy}1��˔�l��)��c��_%)��BŪ��A��� R�O�if8y?�@�{�����i�Q�e,4?VO��8���C���9'5'_�4'-��Y=�+�=�B�������c�KUg�H���3@�0�������?Y-�ҝ����D���J��j�,�w_R�� ����7��oaQ�f=%\��#�Bp� Φ�C�8���
%���u);)
I�H�kA6}*�\2���Ps�uA��#n��W�"^	nI�H�`9$�u��e36T������1��$\���������)�!q,�c�_�����d��M+e���dJx5Y����n�X';+3�'x��I_Ԑ1}���D�#�QB��z��WG* ;�
OZ���b�1hf+�67Q�w��$�]<�L^əG��iIl������l��&�@��;{(�6��ۚ�t�=�4�>�-N�B��J�S���-4M�a�[�$��2�67>�
�-<���N���^ɔD* a�ׁ3y���;��´ѝ?�%n��wp���?��U�f�M�c�Q��B-�5Cv��w+��]]���;���da� �WDloh��x�gy�W�����^߶���wN�dx��I��x�-�E�Fo{����o1#7�GHr�ِ>|�r�I�zyN<��*� H9���9Iu� 63���� #�!)�J��M��:�Q~>�*>DT�����>��!#B���z�:~��H-y����û6m��B����jc
���l׫	��2�.N)ٴ���/g_ x���ޗ��G�a��9�1��f�X�����\�*S�\��|�D�>}N���L��Z��� ��-�~�T|���,1G����W`��/|w��u(�%�U)ю8�Z��do�I����,�rѾ�i-L�[�tQe��M?,�0�I�і�a/a٨,񀣢�V��<؀��R�a@;!���D�;L�飏"H�&͢S6�л8���%�/����C$����"nt
&�X<����[�f�9sB�bM�j��ZBw��2�+�]�Q+������ʻ����{KO�xrآ�T�x`�A9S��ML>荞X��Wщ,L�_t[���k��&:��O��D\���%���{
T�dy9�?'�Զ�u;����О�.;F�!�#�:��ɻ
�l�X��v�u%��q{�hZa�pХZk^�f�yb����.�n@N��K��`��x�%83�Zp�M�P��Z6�j+Ow`�>�P��i��M(%l�I�F���R�6�Z��5v��k*|��R�a���Q
6���_N�!��I4"����I�pN��O0|3�9a��/�1|���|y{=&��ي��e`eұ��~��$2�?�e���v`߄5}H�����P�e0M�j>A���ǌ#lzM=�	���HM�m�����	�}=9�qk<d-��/�b�oӫf-W����Mh�C��i�h��ѳ��?WwB�:h���ŵͷ� �?5�&�#�K9��������m��o�� 0Gj�A�MZR���o�oxm�9.�H��4�2�-�=HY�wZ����zN� ��ӕ�pGd�s��he��_�W���`�FGbt	�H�g�\	�{S�zX7�s��f{�wȵU�:4�]�_`��ؼL����S�Q?�<�r���l�^r��JL����*d���Rq|w�
3Hw�b���Y��	b�O��c����b=��+����}���� �
�nV{0�^K��#��S+�\�1��M�R���1�ξ���G+�Y$$�����\�Q�$���5 K�Q���暞۪q���q��7ݶI&)��$
Pr.��9/L��<��mġ-�Y.�����і /\Ę0\%��#�A�8�Rm�.<���t�m�mg8��Sxc���%r3��!��BμG��|��&�͆7��v��$�}�r(I���"�	�ɹ
:z��[�r��6@RQ������sj	C�އm .	fXd�L?R�9���.��sE�,���\���CFg�ښ�5UG��� {�pY��5�|�+��|G���(%���?f�틐�>׊41�l�A�_'�Ԕ��.�4�}�Q=�C��f9��9v=dd��Z�,I!�Ӊ������N�c�P�d|�4���3�� t����h�7���_v{xB�N��2�(���Ze��z��U�_�#�<�^)�`+�������z��i	���c�F���4���:)��HXQ�M�.H��*�u�*�ߚ�-�O�>:dy�!�B,�("O�%[y��OX�`{�$45�E�T4	4���[�Q$��:r�Lzԗ'y��yu���4�1�,���lQ��8��@�ש�9��4��j�n���E@��C���l�0��)��-=�%]I"�R�pεsR������S�[�f�T���PZ�T��r� c�\�Pr����L�K@��5u�jJS��RI�E�QY)�7��?�� �EM<��L�����[)��V�=�g5N��go��_�"HػS��s=�u{
���pk���E�a�0��q�_!d������Z>�]=w��0�����]M�B�DE�� 	��{��qE8��{?�Vw"ݚ̍g��S��^`�cA�W��*'^�0��;F�7�ku�[�0p�Ù�̓J�޿�����jV+`A��ք�*�Ɔ1�Fd^�ja��yɁ.�<B䅽���1)��˪?)H��yZ���i��vК�||;	YEk ��:��f�]I�A�&�n�o_B/��>��
\���މ:�<�ڣzb�`T�%�sl���U�_����8_"��[���<�^HP��'B,��*�d\��>�] I�E�0�Ur�*Rt�����^���G�-Z�{Jq����A�:G�.�n0R0�z��Oa���?�+���A����30�B��J��!e���W��~�ֶ�vy:;�����/#�u��t$S�'|x�i!]�yTZH&�Cv���y��N6�$�cg2��)�t�gBK}�L�EAڳJ�zS� �R���K8+��!-7��+��ކ����7�7Q��@���AI�M�og��򬗞=�IXbe����kL����o�K��O@o��F�����t���&0�_�����+�i�y���"�_C=1�[��?:�q��6�e�K8�5�{�d��}r�����0��д-.VQ�Hzǉ�KN�E؊&���.�I�3����?<���ӯ�h�2�L�כ�G�GP��/7������^�Vk�E�ˌu
�M�E^)���u��{?�S������Oy�.�U�3���N�bLō/K=��N�;,=S��bhڹ��饘��[H�Ƃ<۹����hXz�����$���I!`�c�w�ob��ǡ+Օ ���Ւ=#mJy��� �OW�>�?sUf}���qշ����[P��~�(�J�@l��iO���8�rn��b
���K$FH�3V���Yv�Л�=��Z�=���̑�Ws3��{a�D�-NZ����CZ �v�Z�K]�Nam|7(T�r���6�Q�s;�l��/�ICYk��Of�l�x˩Y�Uz��+}��BF�Dl<�2W�
�y���w����terG!������e���Љp䖙.�Q�1A��A����4����G����4ؕ�t�0t�PR(V��Wg���I���v�m�V�j����4����^��7�����a�~sGS��؞�����&��� g�|=r?g�h╆���`0+l�!O��Q�'@~Un��Zh�i'��o�VKX*Q?�%��!��~y�pԜH�Y��5Tw�
�h,�d�e�9��+iʅ��Q7�ɩꖝ1�*��9�9��`ι�Y��tU�����l���.����bƇ�@�eV��.gp��|�i�ת�T������*F�#�_�K�9����<��bep�Lq,��R6 %�c�0n�H�pS��LD(�Y�H OkƑT�>0��� 6l�jt�Wwg�%�U=��V-j!�&�����,.��(M6�ؘ&n�*��u�+�,[� b�m@�?O����Pa$S��M�e�E�L�!��{�--3���)ԩ!������$fD���H�8m��K�MEu1�����alP\Ō��<R%Pz|
��!��/�z�7{Bx�WDhY��I��_.���'�t���G�,��S��re�7�s�zt�2����6ܽ�|]9h���}�1�
��=_B_z/տ;J��Es����ʖǭ��(��c)�0�qF�,�%̀��i4C�\�8_�ћy��J%��K����:�K��+/�����޽u�u=��mm�J}?�P/��h��Gb٘��m�.�-�n`.c�Ħ�-̓�ls;l�S;v�h7(HI�I����Sp晰M�(�ph�h�B�����������ٻ �f	�����0"�!e���Y�$؛�%E@�%�&<oۓ�1<y{[-��5��l�V���?n�v"�Z���W�U�h��&��o݄з�k�~�{��e��ab	v��?��]cj\�y#o�G�0�D����	��gZ�cí5��l��%�����Ưm�.R�#8ÏL�}���}�B���9�!T�ӓس���BO#��9�hL��7YxԢ���c^דNf]8���T��l�@�o�A���o�Eѧ��9rȯ��F��� �� CpQ���J<Zd�T��`VL>H�PМ2sc4�X��)]�P#�r�*��ez�D��(s��r�հg�e�?��u��Z.���$?"�;�<�#5'��#f��� "��`�[)��%0k�.�p�(�t��j����K.)�#�� �~��ɒ䪖���p��z~
�ѡ�}R�/EX��˩�������U):'0Pq8��d�=�q�=� ��1ޮd�DX05���:=�V�L�tlٕmpED��֠6�I��k�α��kb%.ɀ|<��m$�ytPEa�Ɗ%��u����h�^���U��d���	�6S*xH�F����7�����mP��9=��2�]G�rtm���ј���ZєE_�7X�[�т&�^�5��k�e��),/q!.
��Hg�}b1c�59��a�h\��׉�.HH[�����8FOt�th�R��|�pD�b܂��M�lT�K`�a(&��7*yB���˽�޷���l��'��:�#h[�Y32o~y�7;����I�}�3E�(���p<Ж�~��PgP(E��f���{W�|�椱KqV���d����Ɲ������3�D5B8p��AE�V/`iʉW'��˥�êl���hS@@u�;Z���	tI;��b$Ɏ×�|�P�B�z�`e��e� �O�DF��.Km�0��4�U�G/I|��0��Lz���)k�13����.�W���nKK��kSS���Y�G�?�O�e�)���_� ׯL��.dΐ."n�rԤ��(�|�6rz$=�3�$�$����4�؏�%���Y�l��	�Z�t+{��x-p29K��3�����.;�e�'l��v���fv�Mg��
C�5%V"HլT'R:ukZ��Z��b�e��ۇk��`b����>���A�����V?g�}��^��S�(�b�a7�?d�n����E��s/f��#h����=��Zb�D�$�<�t���m�7vW�v��1��߹^8E<�*s���c����4�O?��g�A!|P��#���}��ڕ4�������L��d;��1BpQ��z�(�Ӹ=��r�L5�������;��;�Z�J�E\�F��c{�m�L�|�W��[#6e�����tU�"~ew�pZB�*���1��V��"�e�^����ya0���y�^�m<1�L��R�_J�ϕ�9�R{���/�W���q������]G�p̅y�=���|2_����~��n�8��G�h�����O�e_�\��1�U�	UA�2�>���D��GM��9�Z�^����Њ�1��ȸ"�(���	�¥��;��	o��;��Q@��Ί�=u��i�I�NÝQ-�t���|��eO@ �z

h	W�s>�Ѳ�ζ��/w Hђ�Gw��e!�
�l2
�$���RB��Î�9x&6� �� /�y֦�BD�bki$�Y�ȋ-�۰n���9i��Ͱ�<P���+^��A6�����=��}���PZ����9�� ,�� �D��=�E�o�nWJm���$��\���������+:tő�ޢ�AS����� �ͤoca��K�H�Ǜ��Z2��$I��u��'Ѐ�7U�T(�J`�_�Rs�z�3�W�������ڏV@i;�6�%
�XC�E�+Q?������8��L-�/T��t��y����j��Y�g�\�i�,���L�c�2w �����'���u�Rb�Ϟ�mL%��^8c�X��A*���!��D�����a08B�XԂ����r�����Kw'M���	3��A���zWH��j��s�����x!�DM����B�GzQH�B�V�Ă�Q0yg[�!�g�W?��jr�����-����K�x��yC��VɵD K�n�D�A��H0�5��{w��*����ez��Q�_X9�}2�:y¡}�B/���zW?��Ѣ�XIo$3��؃�MYs)�^���K�FW�&ڷ"Sc-�pS����(*�X}�#2Øj`�Е�w��<~�8�Hi���U�۔�}��I��)p���x�������E��!�Or�+���7b�͵U�Ax�����E�c�M�R��;��S�*-�|�uℌS�X!�}��5�����8�ҏ70:|�F���	W>qy��L5���tς���h3S|���9f��&������*��w;*��J�+G!�@�98�4��5�������������:b�1:�X��3J�S�'|���G'��M9;Hd
�ط��
�}i%3	-��c0)4U�U{�l�����pxxq%�!㻎��|;��Qc[��i�Pp�襪���g����3=� ���-��|��j|-�@�93Dd���L�(�F�r���]ci�|�E�ʂ"�Z&���h��6=K�X��#qՌG��}~oS�i�^ȃ|I��u!_�5�S�����{�*!�M���y.`2P}����J����q����H'd1UM���22V%�:����7e��cq�T&�r~c+�6�*���Zz`��d�]B,��]������lo��<5W^�}Snes��5�m��k̘s:L�W(� o��xu��3����͆\`�\�C"�0$�jr$��]}v��ϡ?�\<^���?�����mػk�C<���Z-f��Hb���prx��9�»���3U֌F���ߦPi+6@K7&dv��Y�v��Ť���{����OHu�zzv\�\��x23���_��V�QUsw;5�W����%=���&TC�vs:���(���-��̠Z��	�/���f��c=��-VU�D:�^�N,�rqu,e3�O@C������*:6�o&B��r�jKӿ���^8ჳ��q������:�F��P? Q�� s�2�˭��X^��`���n�/'�eꈕ@'��T&۬�Х.Y����l��jmUi|�]%o	������R�C_xH�,NJ�V5���}�mK�7����087i�(�X�G�Dm����ub�����:0c��'l�� #kZHτ�Sa�z{gC^�J㪓�)@���ּ��{��^��j� k�n�n1�Jj��u^X� x�Nk;�Ec����E����.1.�V���d)��>���@|�?�W�X�Iɐ�+����j�Us��E5��>��tT��+.h��o���}	i ,�<�r�S� u]Ծ;�٣����Q���	�܉f�.'�e�g.�b�U��Hh�������k,��՛�sO)r�	���5Y�/I:Jh�<�e�L�MG�Ԫ�f�+j�B��"9�c=!"����� �f�*��g� m㤒���%4�J�^k�៾^���VfB�ͱ`�y,Lh氕{����i�g��Ώ�]�,^�IaF ��|�����E"��1���#0>I^����n�8����#ĈeNE��|�L���f��(������2��)0_\C5���V��$6���&w�>���9�(W��P��p�oQ��=���M%�.����b\佳fٝ]�&|G�բ�Ǹ�Y ���wA��]x�R͝��+��"��D�H��U��HR�w�2M�U�_�i�,�uO=r��� ����պ���	P���EA�]j宒�v�����ٯ�1MTD���d!�H�L~4����(3��xW��>'�zx�ㅳp���ơ.��-�	�K��4\�
�h�)�2�~��h�R3K\J�O0��"Q���=�o���v�>p�R|�I�_�y��U��♧�μN�aL�g6���~E����ɵC�=u`�Q�'vvt�$D:��u��ǑCM�B�7=$�x�ӑɘ�2��T�vu",B�SFD�Db�&��SO:QZ7׏$���I���>�NQ̶{��+���j�ē�vڛI�
'�c ������x�orNSѝ�Z��;Nli%XZ6�{�&���|XȰ��:��l\X���?�@/5T��c"���K:�����p&�Z���(�"�c��ưz^X��yN�`��zp�m� �6�>��e���3����]3z^���L��	���oWKx�?�3)���ڧf�~�(G��c��Fv�Z����}8y}���N��n�1����e�����e�z����F��M�W���v��Zx�#�?��k��C�D|���B
8*`�[���qt�{��
���&����I�.UV5��W����l��,py�	����X
��B2��@'�uӗ���o l��U����J�.�/�cl^��/	bˍmW��K�֐Ю�����S�ar!��k��;�TF��Q�
�����B��{���[���^KK���[�i��N������9����Um�v��>迬/u-����o�ON_+�j����ή��W�P����D��c�V�O�z�HI���x����H�a5UP��S��ћow���"�����>� �?��陮tˮ#�:ϳ��{����"Εf�z�A�y�=>��{����^����l����:�����ɼى���t�<k���če�ҭ��Ó�B��&m�ŧ��κ�\s
�V� ������6�=�j�>�4���?�D󟓲t�(9��Jի;~!I<�>��_���sv�0N��,T`�~�n���<T�hZ	���*��<c�e��#����߭.Wͩ�M�/�J�p ���|RZB �-Ց��ܡ�u�_��M����1�C�����1�M�'P!V]�[�7��<�P����`Fx b�j.s �>)�讎DL?v	��R)&m+4�Y�h��1�ֆ�ͣ"oi���j��^VOݢp��7�?yԦPޗΛ�d�� ,g��o����CA��߆(����j�S��Sߒ��*_}!��E��� ~�,�"��8��hl�є�`Vy��0/Mp�Ga��a�[�P�;�V��x�İX�|�>S�	;yID�녹��S6�\����iC�����t��ڵ�l�w������|dtAn1��f�,Ѐ��6��4QIm"lŐ��2���7)��O�_f2�bЊ��J�Y���$�Z�t�������S�J��2��<a ���p.��dé��u�M�C� ω��k���O�����ط.bKoo��R�f7DMaS�� }��ז�XB釚�Lо��	�R�z������m�E�"��E�AX�_��,z%��E�G����i�BF�P�>V�����"�ح-��@�?W���/�xhmћ����%��ov� {�A���D��!Q�/Z}�"q���[smp��O�D��]�b%c6,��#����dl�iG��Z�=�*ǥͻ@� ��3!�ZӾN�<ZM����~���r3}%&��S����%?��UgǢ��P��j,��R���~�������䪳F���#�}��t��-n��<?~�Q�i81�R�%�`\��ꃷ�'��tF�u�z����^��A��.�OG�J�:7#9�����+`��G U���r���/-����n�@g�f�^��p�E�	���ڎ�Rt>�6��,��"Y-䅶�Z�����m�2�|9�n{��u?{;Gʤq���x�}֪X�����8�2E��C-��3=HtsSZ��eK�W���ф��ڞ�:I�/Hŭ"3����ʬ*m�i92/I�d���${��T+��~f�������& 1VUݱuk}mT.a��]�Nva��ڈ�"�܃"�v��Ԝ�C�z�M0��Z��j�}�\<�ͨ�(�C�&hs	����7�r�ڊB�S��G�[܁H��>�C=�S=/�����P�vO��{i�o��]x�iŬP瓊�:�6Kay���)��!Xr����DK�N�L���\ZI���\����I어�6� ����=�bu8r�Gl�Ư�/7$�H�̞�o8VY���z�AVu���T	`�e�~�ЧF���5�a�
	x��3�T�$�����=	޲&��@ƺ�\�*��<�I���YO����;&����l�;�XB
E1 �l��1oP�ߙ^�A,�����IdY���� ���}-��z����z|ӛ4���8w����������ٔ�a�[Z*���u@��s�w#�p��&�=c�{��.�s� ���������L���0�&l������\��w�u,�̌<*u�@���[�*�V�H��Žj��|���L�����*ˣkA��o��9�T�h�{}������K(��b_	�!��{Fb� �p;��3dn/����cMCA�a�<����P�'�Y�/8<��ȼU�������8�̙���Ky͡�v|:$/��c�l%j���X'�YlZ�����{�K���5�]86I�?�J�I�."eӫ�Y��[Ɯ�%&��U�n���(l�<o����K������ED��pY�}��WС�^�~D��Z�A�Mϗ�G ��wzos�o_=��4!?m��>S�И��Q�2gs�C��]z ,��L:����&��MW�R�UQ�;� G�,HB��3�q��^�<�p�-"f@MFNy��c��1*2��b�w�a=56hӷB�fNL!#޺ʮ)��3���}u���6�.(22��z�4繈//���p�Q�;��O`�vcd��0���y�{�nf�䝩{�m��Ä]C@�K���{�������B��m��������`H��sN]	n��P�';s��h���O8��%�!��B{���)��J�D��&����D:���Ĩ�.��h�h��-�e�a�7V���ε
8��KX�M���Tp2�:��.���312|)x��!)���}$�8����AVDf�P�BS��.wpJ����ǧ-����5a:�	�Ix�����C%��G�A�$�Վ0F��Ā��`�+%g��g�ۘ��Lj����ڬ'�2��0R�����n�ȑ_#x��8�8�q˯xuS��b��j���l�ʁh � �@���Tn��1j;����ɒ�U*3)!�i	ǂ; �o����?�xo9�'�T�/�u��4 ���>M}䄱D����+�c|�#����9s���쓷I��*���!��R=��lI����������<�v� ;�y�!/ZF�%u��e�-�6�����y_ܓb��b'��\�f����[��������P)�Dd��L%f{O�uX��n%F����9n�P(+�<��s�;%��k<�ٖ�.ra�l��G��\Y��w�Z+���R
1�(ԛ�}I��Lu�g�Jnf��c&>�>�N֖{��SJ�$o���A�Y7A�d�9iz��Tl)��Ρ]�'�+Ŕ�F�E�0�b+f����	8�g�A�`Fr�����Di�?ݪ�9U�d��y�����u�V��M�]��v
_�I�"���׍������m����*
in�=�%a/H��8_��	�)�pb���)�/�p��Y�Ӻ�>�'%��Z@[k�ϼ�2;&}�{hZ�hJ�U[{� ��
�d����'�vͥ<
���93|=�	f?�sz�?���c��6A�}�q]:l0����0��7`ı����z�EgK�dU[�"���f�@Vj]��Z��!����pIf��$��hysY���GM�M��$�"��\��9G�Hh�Ue�xt�$����>-s�d��3��V!_��U���U�txtb��2D����L��u�ғ,�Yb{�X,�x���+9�Y6�!���0��nN�0�Wҵ�[���0�:h�"^���{-4��@Y1�9S���G���d�8�t�M�o2��N�d>��#d<.���b��=�Z�}�+��q��NOM�-.=}d�O&��\����kw�+���������E��e�xB}_Hܖ=��)q��U���f��}��.��������@����]�!7�N�w��Չ���V;D��ne�N��3��$s��nF�5ʪ���H� 4��f�Ƹ<��E�6�֬����j�OE��T�t�/�h.�Cw\�^z1��>X��5������9�y��z%��ZsA��V�/�L�IT��=ؑ_j�s�fk�>��1��!���8#�3��T��Y�;̼Q�� �w���Ϗ�R���!w�!L�T�B��@I[=�ͨ�87�DiO����A�����gXIM�|�ӝ�.�O�T~֜���o�F
ĵj@�C�U�_8d��3�J�T��ܔAC7�m��+}�U�ɪЭ`]�e" �s�I&o�~�,�I���+��#�k)/Fܨ3=��#�-���ޤَ*o��=��v�n����[���(�U������2v���.�ek�n�=k��3Bkyk��PNRI
=�p��Q��8����Zm'����_3r��m�v�f*�.� ;�+��I�;kI8�[����c93����6����]���m����9`b!s]�/�������ߘ��?vv���Pw*52���;��o
Ԡ��e�B>�DJ\�{�.�$��{l ���h�40�N�O����G-ً읧	��PF[��y��`#y��E:��ղ����N_d!e�w8�fCb�ڞ�~g�ߨ����m,��k���G��>T)���;�hb�z���wG�/�栉5hn[�u���[px8����8���L��uT�p��[o��ԧ}�Ӎ�I�Q5H4h�Y���V���\z����j��C �G�s�}ц4��N&}�(��k
���_q��
M���I�����r��CRXD븨k�Ug��ޜ�[�	$я���-{(b����F���Ui�SF�A�kbno�uz�\�9�Tg��V�??b�d��7��^.3���k[f�
x���j�������B�Jl�5���5���;B���_��/�")��Ji��^ ��X����p�X�����Ѥ�i'�h��(�� 56R��KTB���V��Uı���o�I"z�#2�=}*�u�#�G@�\^��8ڰ6��ȅ�� �9v�` ��^��?�$eo���s0�r"ʃiU'���3��L�-t#��Un 6�1�<W��N)K�Q�F��Ց�1+��8�-v%<�9�������JI��d���i�9�`�fi�ǋr��|*�tHi���HM�C�W���q��Ĭ�)`�&�ۈ����q#���E�E�U�l٭t�e:�֋���nG�N�2�S-��ܲþB.�9L�	
��mi�1�uD���?SN�<ٿ�f?��]W�F����폈�3��~� �س��l��+h�v�2�*Tә�(�
G��9�,2��PpX���u��h`i�Wׅ`o.�9oK{ۻR�n/̜S�/�ĐՒW�~�9�=y�I�[�n�$l�}ǲ�(��(�+����V*U�Q�oĭj�j��v=���Y�ZF2�
�Q�zS�$�9,j��{N��=g��j�4���6���p��'���[���*y1N�	��ދ��L�K����+��ӟ�<��GO��D�
>����Mc=���'�ѩFFOpzؽzw�����{�/��)�#�{�oS_�Y��ky�%�k@�DD���X�Q����/��T �`A�2��c�*���w�D��,%�<��\�K>8/�Px��� ��d��5TRu����?y��̯��d)�.����Us��L#�A��٬�)շ��u�R˻P�������~3:��"�/!�l���yc�h�p��r>~0��pq���m�*B�uk�Z*c�%o�C6fv�K��uT/R߃���)��M��~
9���GD�c�6��������R�������9��H'ÈlDa���7=�|�"|B&R��)��:�]"ܐg��0�k� z���͐)O/ԁ�Q
��!Lj�b]#s��~�����1\��2`��1#���+J2�� ٔ9Bmj��;�Se���"V��9c�͏�Y�]��;r+�X(�y]ிHWt��d�xS/%�vg��¶�e)�AG��j���gN�x�u���V�-�MH����*4);2�Vǋ�0�NQ�Ɯ�<�%�t�����M̅�:���)�&�q&P.�a�7���N��^5	��I�c�U���ģ%�m�=�@�',�h�#��R�-S��j~��&VY�Ԛ5�̾G��8?�-��!s��8\o|�t����p�?N?1ى.���"�'"̌xuF��%L稟5� ��᝱f�0�p��e���tc��؄G�=���xH��hwk$�� ~��tS:2�L
�/+��V�T��P}�Q׊��u���7 ��cf�'^*:�"p�p�\�?�}�R��jaX�7����2�H��3��,_᳛j���ڤ}5`�ؼ��S��J���9�M�I8ρ�C-#]N�a��)s��䇇aнzX>�Z�o}ȣ����ѿ���#JuD�F-.l4Q��]=W����=�yM�� v.t�]p�-�?�wis��/��Ҧ��9�S�l�K���2QFp��^B�Me�1��U<:��wP:�2ú�+YQ'8�D�11khԔO"��
���}*�)��0�6�*�KzH�S<��߃�3tt��N��bס ��O�����Q���L(��C<��������E��T?��bi��>�Z�f�;g`_в�0��f�à���f�Q�c�y�#{� Q+�b/z����ngt��|����,��8��7�gT�'�kUP
�[�׽̶E�)�o&�;��+�ol��r���Rr�?ͮ2Bf�!*�����K'��퇅�C��T6���0�F�k��)�p����"�+ɵ~XK�dȹy0�T��h�H�>|9j�z����|7~����,M	�{:}�揵�U�UA��z��IȯHXrc�Y�yӴ��S�|om�f��V�Z!54�� s`�V�:l'��u��MJK���%��ܠ������(����wz��(H��a����_̎��#���H�s�gx]L�
����߈����(�8��;t��߯��."V���5x{q�������69jߛ�GH-�YrI�ǭ��73��[2t���j�!�x�~�H�I����vKE�*������_d��y�����?���r��1T4]z/�ǱJ6�煮�(1�PX��T8t .RRH�s#�Zn�[x��y1<5�Xrl8!��*�ys��� �p[��W����2]�a?�D���A#X�w��~L~�d&��T*��O��z�9ʇ��!g�(����0�E�~����q��t�Ì���#����Vh@ �� ��_���A|��]l`�O�u�Y����`��Х,�h�t\��J#H�/�.m�<��uv7k范S-��q�b����Ez��!�T�kJ�ߌ�T vM�B� �cŽD@��-y�@�ژ�q��N.��V�P�#�Q/�����6H D���M�kY���w��1����EFL�`��ⴇ��1�p:3=�wI�E~���H���D��́ts��^��3�&bC�� ZL�?��5`�؄�P 	�Vj�GI��*�@�"�4JE�M|M���^�߿�:�o(5��~���,+��c:�� �DZ�Uf��ϻh�`�j�
�[��)^_#k4�M���Ob<�/����dܫmpr���哻�t��D�Θ6(=� �m �q�ŗ��t�n���"\"�b9��\�^�,Gno����j�`����D\2t��9�vQ�����V���#Nќ:�}�u�����ǹmݬ�U�*��q�O.�(�/���(I��9�q��^G3=dc}A9 �9�n��l�2 ���-�t᱌$`N���i�5@X�!zsA*YO�<�e����FV�mw;+h�cx�_{������&��͒r@]"a�n��������4����k!j�>���-Bۄ��a%���� YX޽s��W�p�{%���E�J㼵(Pp���
��t XP��d��Q��iJ�8*�C��j�Ze���WJ%����xwvG�[���,Q��V<�?�e�M�MYl�ċԶ`�â�\{'	>�g���U�ܬ�����wDV��M.�˦#Pt���y���&?p�1��G$��k�4���wW"�u���{O�H@5jJ���*�r��g:���%o.JG�%4��:��A������+I����I�[� ��{~*wL{�9`�a"�e |�aA0hO�g'�� t�A�N2,&2秭�g)�>���X23��y"��H��y��������LR�oyV�$���;�����c����2u>�����kN~�_�-`Gl�b�uc����:>i��G�� e�|�Ksq��[?�f�6�����2���^M�ﾸ���8r�N��	����u�K�ɡ�iVN��0��c�K����pt��l���@
E���)M�-Md��G=�Y�Rnn����������BK�FM�Q+�С;âH5(���!��8��r���W�n��^�'Ff��Y0�<WJL	�q+��"L�����bD��^6��;��(Ŀ}+6��W;J��WQߔ�[?�9+�j��S��V�$1/��W�ȷC� ���M���<�.ݫ$�{��	Ȍ19�95�C��o�c����3o	~Vﻖ�p�4xQ��hոKD��R:���M�^!9RP�'��M��,UF������g�2�DW7�j�vD@�аN1�X��ߊ
��L�p\d�YȿP�e�����	H�o9T&�l�9��x���Wp����)tOVe��~�{.�
���7��Uf=�=$[�z����ϡ�+�'��{�.Żj����e}V���FV���a�y�GM��l�����SS����N���7���E��o2��SL��DP1�{�	�!2�����o������lHXi��x��lݞ��[N���c2����nâO}xmd^�����(���dqȿ��Kq?7�W�֔��_վA�q�G�=���,Վ!��)s(O����m�["�[i���r���"�gd�����_F��U��B�C;ssʴ��8Z;g��s?�)S�L����!�t��}���Z_���FvE� ��pL���FL $�kQ�1w�K�[r*Yf^�*��d�A�����sa+4�!I[W���i#���d�/�R�E�ڵ�~�*q�~� d�Թ��82O�.�Z���;��x�%�U�|C��~u�lWSGE�M��U���mX��C)��;�PpFW<xe�����Z9���A�ѿ�����}'��Fh/���$�/�"����HVe�2r����M��0
�-�iM��
o`[k\�d��)�����v~г�U�E��I[����2@(�{(��0 �Ϩ�?�OK���/�,`Pc��.�o{�7���U�A� �w��b���My"V^Y��/�Ek��*c�m�d?�@��&�y�������2��?����5��xM�q�S�/~f��iK���)��rڙ�l�2���3U�E,"b��<(������}N��Q�@y��f^�P�Թ)��z{պ����l��u~����$'0Q��T�r�m���>�4uY�k;����G��x�7 n�-�n���ћ���B�������� �h�2�������$�>x�n;Oe�	��v�q�jP�tO3H8.�G�}�||{W�����������`�[���<���5�V�u�
���{�ŜU�@fY�>�#*F��7����&AO�?KPk�5"��Gl�P�_�b��b�=�����]Yړ��ߨ!��!g�FJ�WS ���]�E���k�sz���@�i}
�Ywxﶺa�2]	�w�����r�&	\�]�Y��fR�̿�@�5R2	.qհ8�R������'ǧ��ȋ��PD��a�O�ʴ�ؓ7?���d­�#���f� ~Qyh��M!`����R��`4sZ��Ew�'�td�)��7���� 3~po{m u�̋m���F�j�}*WC�2�x�"��Eچ��������l��$1.��$��	U�e��B�+:-3�IL ֕92�l���#����_k~;}?�K��$�Q8��KI-���GsO6�G�鳦L���;�?$Ӱ��dU�i�T�eOAsP�rO$'�+��
�`�<������@��B~�!��N�b0�*эX�R������/�]�k��)z�p����Ď\�g�׬�Փ��)rZ H���ZzF�z�^��(���6����(�V�Lkm��u1j��F��`[%�OS+�t��M��h
RjW�_j �q�y�DR��#�����ghe) + �c�A࣬�KQW
��Q��={<�<���7։H&,@����V�m����a��M�z�Ueֹ>��s��[Э8�B@o��ޮ����V�y����LiTЭ�W4���DܦbVm����zU��Yh�(��i���\��6}V��茿u$��HT�b-}���8ŵVYt�%+�kc��?����F삧��M��C�;��|���3�[��&�D'�3OzTZ���	��l���q����&��۽4<�<��t�YW�R�~���B��3�~ןl���Y� ���b�1�7�c�ݡΤ�8���c��&bE��}�t�ֆ�`���Q|mg�K�e~�\��ޏ*�@��%L�	��L{�Db��v3�뾼��*�J>�%�IA��PD*|]Q4��h��ʣP�· �8�FBN��~#Q�����7ӌ�c�[�-��C#ߝgߓ��1�_E� +L�\�lD�znKK��&W���4�@�h�}���t
�fItY�`m��^S,i���FfR�$B�­�b�0X]��1�*K�wrdZ̨=�m_ [���rߺRL��8�h6o3�y;bǣNʋCl(�w���%q������x���,F�2q�e1.�"L������b�կ��A��+�^�e��f?�'<#D
e�.�`�-o6��:�Fcz݊?b.�h�$Z��cT�ph-%Ņա��͟[�/��:�g�b��";�1ȅcSC{l
 �oHj4��ڑ��^�[w>u�`�E�C�aaʙa�2�w�R�@�芦�Y�o2�Ҏ��? ��p^��cVen����lКo�ʨ�6ɰCý`&yN�/�	©�����m[3u�t�X��֦�P��T[1�1��k� FKq?4�@��ymv���侎��Ԟ�[�6i�&dT��0]>��ʄ�Hi�f[w��'���p�����l)K��h�Q�ч������{%޹����k�QU �����M ��Y�ɿ����B�h9>̆�)X�����S���S]<�sf�1'�<ox�z�C�z������;�Hϴ�9�2�� bI&���y8#��A.Gߔp{dJ�DA��	�o�n�����NO��+f_|�iJ�E̯�x��e������O&B
��IzC`/p;=/���b��PL� ��Y�Vn��q+�ns�P�\�I�P��u* 	��M,"5�Uj2{-o�aا��(���*���V\�,�H ѕ���P�La���p�����A�2 
 q��|�D�۝�](��/M�C�/�5��Zj�%��$��U�'��vD�hY�bv֖��p4�PКb(���<W`k-HЕ�\��f72�D/�R�{����oG\@m�FƛƃY؈y�֨�vD�ոX�q��aS�� ��?yL��e�D�����ʡ�{�n���"}�T�ݾW
P�y32��"��Z6H�p�*Ũ���|���]-�u����� ���D|��D��]67�����}:^����~�����2���K.�uWl�������è�D��wEe����b��K�+pRmdzd������3�A�s@�� �r�q��7�̦InM#o}o:�
����*��5?a� Mp�t��lˬ��c����	C�Be���T��ƈ�1��7�|U�Qx��ՎA.�)�5Wt9y��7/�Fzx2v	@d��U������\i���F:��\�
o�k�����R :���k�4)�����zM,F�$������}~�Ӊ�R���ڧ����3C�z�nn���^�wA�����df)��J�c�~��Kk����t/��r��ӿT�$�״�繡M�sǣ��o?�<��	���>�3�>��%1,
J�]�$��K�P
)j2x�����m���?����[�X�D�1�����Y>U3y��L�_c z�!Dv��-��-<+�\(ܰO'�>�jz}Q���|ׯaG��C}��}�-p�7!E�5��4�N��Nq�y�&����F��$���":�KwCB��͉z�ܼx�H�U�?�_��Ǥ�eRN��E����9��aT8��s�3�VS�@f���E� �t�sgZtZO�
�ꅙ*WnO��s���;|�h�͛�(*�8���9$���=��;<����x�Hvi-4�Ȳ+�Vv��2V�(�{����0�8�b�z�7(��v{%�Ƥ;�f��C\�"g!�&Ө6�
���R!��A���\<� J��op&-������N��,�Js�V��^����]��jw��	�<���n�jQ�M>U�d	����O�c!��{��I*>��ؙ��I�[U����hh�R�e�&�m ju�X�v�Ȇ/�<��w���`M�.kpJf�4Vl�AV�@ 0f�zd��UH��j��&���*
_#B:Y�x�/i���Pƙ'܋r P8�YM����!!ĴI�c*�y�֡U.+0����l��}�Nڈ�&�"|ٕBT<�3��^Z?R7H���&�)	QvH��_��0Z������[X$C�D�ms2q	���4k��ƃ9��Re�.��R����̋���Up�Nv�D�Z�;����UW���� $�������zW��;���k��j��(!)Uw���8�m�3ݤ/⾧M�B���ܘ�/A�� $A�H�����kҽ��4���;��.�G0����Na��o:��@)j��n;ф(h~K�_����D����;��f�����H櫖�w�Ñ	S�:�g�q�Cv5�>�3�F��Sp�7I�r��S�,jp��GG"U���l���"����>wƑ_�'�1(�XOi*lR�lM���PH����N�@E�J�n�3�#z�t���~2�:��J��.)p����!L��&ݪ��|f�Q���"\��� KwC�W��^������ߔ��M�����
�3���;��z)��#Q�?���)oY����N=lpY �W�H+ L�[A
	�4ө�za��ل�_9>&(B�����lu�9������:oɋx)f[��=싣#�P�[��Ez��="��b0�3�>K	=;x�i���9�oi�jEsO:�,�C��M�z�W!��ga������>���)�n5`{%h�f�#���!r`�g���W��4T1�(�D�U���zd�z�ȅLS����N�Q�C?�q�F��CJ|d9A�:�hW�㍙�
D�����E�}��	�f1<,���c(���b;�`U���4������w����}BB�\lN�ԢO@V2��$gnX+5'Ǵq���C���p���b���>.M��r