// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C7hPYzIQF8tCpvWhptpkssK+Ua2GWWFYxG+RzB4Ym7oxXHMsCvSvD4m5namVMaIK
grx1lbXi8q9ITYQ4GjchIn7Ttd54mhGho/MJKvrxN8o85q320v8HIzGTwE/AHxOl
zsPwUlu0HoTXA835bHxt6npxmkQ5LfbTRlpnQqqIq1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
O53X22FbLrwPEZwKdtiXvIafLDpYsMajUmY60wtF8GAOTXwf2VMdBwPY8VJP6eO0
Nx3Pj8jxbC6p46oTACQu8evVFaOQiGq+ZoOEGb9PMbQoLa36xHktWwyUFxA0tcBK
4jhhO9wgwY3/HugVomHQzNyW6odvrbh0Rd6lbNEVTGYldx4+7xFhdVmlWKfluGYz
74oA9Ic6LnBiJ97tanvpQCp8URV/0CH/Xi60CxUFZkkTD+OFEquiHZkSrN0wRj19
HuHN2yJLY8a7kphsX0GS+GnQCyR1W3r0111le5yt73XgBoT6kmgjPanbSUVT/0MO
JSsCelxBgHb7HBfEoUZlWWWOckcV9a7S6D1x9RJFPpBPxSglj81Xrg7LOkts6oko
ta7dfIVHtPFiW0vSzUOq8CpxhYJrlHO7mRR33gqRbKTtr9qF5lreTO12D6//l1zK
2w/o+0zYRxlJEdSB6f7VGgncySpkwe1lgXetJxm4Ck9sdXrCDKCh2+e+AzgNnXu6
GD+D2E5YXMbAWFm/TWFx9vCPVRT84tO43i4L6WvcZFFvzCXk6+uZlBa+jkF0MfyH
LjnoD2FMQli/0XHzs7ODieWtUc4Ioh99avFB5wn3xqNeD7gj1SELcB23waFZLA+F
oXbM6wf//b6rptbzPAiq0838tF2ccxflbSndYY5gizww49PDdgbhkylqO9F6Fgw8
jJgaHuaxeiTLxnvxMyInO10tOYx8D6h0+bwOoDEp3rkF7udufDDu12IPx9ImI7LW
5YMR6mK1KDfbQoj+Jo3BNXYTp4C1ICjJxn3i9gzO65GZN0NkJRvrD+gy/eR9LNHb
9YdW7JvwCeVcYyUbKn47l+sWmLYplCE29gUkKvVnmccWNOf3Dk7pv5JZ4ZWHZF59
1W/ZWMdllgJOyFKjKJ/UPjbszEKn6oT+9Zavt4Xq+POWcBqHNi0RjIl/gFs/00VA
z6ikYc2ph5lpoY6Ak6U++Vm/0QUa2A4BiOPwRKm51+mNaoEVb9W8vYoN28aRmWAN
2XhqkolN4121N0C3vfUujGsBAyB/NmBlEFO9cVxsRQDsO13Vd9N1xjnxUrkQFtbw
agj8/eR1sD/gz72wKbcjEPYa+VOCriBq/XRjkycWeFDDkvLtjoT/zncdYuEbQ/Et
n3jakpQmqRiZLYbHS9PyAsXYQ+XalBYMjTAGrC466aP7Zx3cd29951Pb+UmuZcpE
uJuxdFVcBfctpP1WWxWrfpEaZsAYbBRMLiclOgMsiEgggreW0I7yqyE1/K79pP/x
vlZc8w/Yf7iVX61SJ4p2Owd9jEhCohO4xKp4VEez4zYBGe+BBf2Y+/zSffNFrugh
I8+oWPpdyVi62jwPQkw8mobBvs792nSmgjmTX6tmkjs5uRZkNu+D72qYaoImg15E
P00RkFEkzzznTJC9DLL40fUS7tLjRAl31E7YoKrtk3ELmCSTOvtIduGHe1HIiPZs
PHEIKgTHaBD/S7Mm8dPKibK5tscpaxwv4FZAy5SMVBs/5/nCjjNC/rtRFi6pxowj
7GvuDSiQBKARTC6v0gqwFxCBttiZdIxfvW6Mwjnz1fSxFlmTYND5q9SULnCjLhMT
rNuvsBxOKEH+IXc2XOjsN3WMdZcbYpSGOXd2yXzm7nLx9gsnI3o5rgFgpi1Su43G
P6TmlE/ujIh/K/pdunNHUki7lgIOhoLUsU6tFp/8oeP9rqlMM/lBAQy7rZMY0jkP
H0W8dD+TgujBrW3HKctZWYjv/t1w4nIofltB+WRDf+dUwAJ4wXY8+pJa8fokCMyL
2FACNTFp9LIgWW2Z9cOFxQQYgawsSKJmS/Y4We+sjanWUXYCwpZ+9tR5obmptMUI
PkweDBN2f8hTGHOSMocKu6wPSSJz+xN2yQiYHO4pvhyNwylrJ/9lfv0Wx4rQ0N90
Cht49AsuJHV34zkAbelwu8IYcK50suc3KtcXrBOvIseeWcWU92YerStEFXqz4VY8
s6vuVEferkl4W7qB/fmQVIWfNQYdO5KL8kzoqTxkBvgZyPlNaZgWbMBcLxk0rmX3
WNRAsxsyp4/8q7KytyNnrOy5s8231zzC1maf4ltaciJny+qXmD5FRkW4YokkSVqf
LVduCgF6lPlcjGMnPux7eSgccSIPwAiK4UL8y8uPEDbHrD1l06Wv11T8vczQbefi
cpjCuwuQSMuZ/eT9STXOf9w7KkeZu3l0mkOKzU7ArGvBF7/qg24fzVPqpDIBfoKU
+wUo6uW3yVCY04SQeQml8Dx9zGueeP5ERYin/b5yrZRRb8fRn8mPamO8r0t9D4Q1
POnqCLluBABwNBvz6WHrvdoUBznSNrdH8BnP5SUZ6SoG5s3Sz2BC8xTjHDHvy0YH
eKM7nHIPFkEFErwbu/NVkWRAVHqkKf6I/VW10rIwSeAF0uLVz8LnBnx2X5Or4cs/
RftN6Z9gaT09OC4NJ9lf1ihg6vglqusAmkUDogcQX75fY+aK//IM1bcGeZ3qzktn
7M9Jp8nmXmEw4zLIT2XCLbomugtPMTNpHll6pVNuNnjM3p1ES6bxmyZvdW8sgBzQ
fAt/muMxt0jRpt5Qxc8Brm4n60uVz4SmY7FZdZQUwn2FEgDk5Bra/Ub1EQ97S31a
gWMJTYFwPZgIlPOPPSgjbva/9HJssFa9jdxmZReB6IX51gedbP4ap+e11NgvZCUR
DpLp5FJkKyGVas9b4WvSxka1mkDewVtxu4WOeRKCCTcEgdAS9Qu6Xxg5qIiBkOL5
qGngHmufj2V11HeG9yjMA95/K38ZM5xIUnig3rQoAvFOumFTYZ0kKwIssYLK9yKE
K4Hu5L1OONXBWQcq0LYFls3qlz7w7nCVQIS2Eh+CgclzH1JUi31nEya+/xhNC+us
VgNh45siXODisgV+1ZbuTmkD4xx6Jjltp/SYaxnvSiOGIydts1YStXsGyfBP4yZP
23lKx4MdUeQWHWXLIeYrK3WiwXFiJU6rsyisp5s5Qy9zwklf8R+WWFNe9rZBBd6Y
YlDnrgTWUQqf07B9dchtC8fQh9jHytkAwi5x/kSHlwunBWzxDXd/La/Q9UO5t+b2
uKpYYkw7PPlNILS6GzC38vns9hs96z8h2dEwe2TBmImbDD5UZbKO4KLvSm+lrH8q
Ff3G8ESsiXuCKok82ip9gkdjiLIf5hNqkp5NnIyyncr4TM8g17fQQuiXK1y2AUUh
4PRB7PWN2cEysuSyIrN2zBtYMDVWym+sHgtzCj7JDbUwJBwnUKh9EJsSZay1S+LW
ADh1fnCB1uo5BLvtW+7uppOfXRAqa0W1z55TQPiwCmKntYZxLb7blpdDda/eM9zC
XEo7ZEvPan4+NfLHbOxYYVyg61jTl3T1Cd4MkWROTk0SrISeOv5oy1rGUuVsAqTa
RWJQtPlDlhBT3rIGuNIEURqX6dWxJ0kzllA5fA+UCoG+q93FKJniCxzb74Gj75ev
3ZF9J+JjkKZE09QYvGTDyWPtprgbf7NvWW/38PWliIUthzJs8RzWb7CX4YmNEXyP
hWZr8Y/QjaxUBbSMGwjBC2Uz5nB8HUBjBtIzcw27ctcj8qwoWQ11zmIdl5pUkC2L
YvSqAuc3/dQ3sIo+P44YcQ/ak1JGQukExZeNWy7KhdJUx/UcKFSPruJBnFoeVG6i
BJius4wTuoG042qzH3bRxTu5qFYEyLZkYKEOy7F0N85es26hiwRTEbVOP2FfsCxH
yrAkGqjnjWXNDJrRrOd6MQ3mrRUzpVLhrRdm0Qx+1Po/s6ZBveaijT/aLhU4CwM1
5weaX3VproWAdB2HlTA0/Z/Jyya3JparcDIXVc62u6myKWSS9Gk1SCLWXFSsGwOo
TzpWIaK6n4P6jQKggppxO4PX+l551vMV/95UTr0A+C1ZVlT81G36oL3Y2JK2j3eF
466Jney5pXiklXo0dJtLKrTGu+lC0rniWLP3DJ5SNtBHr6+zz7FKd8+DpL+74Ywj
/H/FIrZiDjMs3YObhspT6b9VGez7vQTc5RSLNZJxUEoYjKmivqhMkmXRBfU3XU27
mGlUTEOSefTM74IjJJb40J0iHeopsGUrT19dYVpFTrwJCELrVTiejttzNfoyQUHO
Flfd5FLp92/qnU8QuEk0RBgHKybvgMos+kQEv6YuZNebSEH9p6Zzld5hCd/3AjDq
27eYZLQZBFl3QuAIEUqrXx7zsp9JWO+R8TlFl+AsGpNRUTIExYnp1TBhlZHnBic6
b2uWS4URDUuiCAiqIMnVS95VFQRdoTSp7P8pMQA/V4DzHG9m9yBXwZ31g8R7HP7V
MHiB2Ew5iB8Grr54nr2S9Kd6Yzs7S31bDyl24DCLuqev0Q6J0lL39ShyUXJgCxNk
9Ug63GfZie0zkYg7lAuVb3r58IdrFu8Ydmp3pLYlvl76cZFidLxJEHGy7JjqcDqk
0I7svXzfIo/sc8CNPXnQIlaGFsNgnxC92W8R7hHTC0fchpk8eO72MH60+FQN1VvP
4XGpAw/QP2SAgCZUjA9OFZMmfaTr2My84C0V7M6VflWNgGP/rRz2MgQG2ofYcLJU
WgOAgMAnczAXdeAzfRgtmqPONYjgCUiz4d/0oGZEEbV9ohBuUsGPZUgCTneED2EX
J67AO+nRyEf+nVyqu39z+KLMEXr++6OIRxU6CCz22Ghbrv4Finuv4/yDxJqIXikZ
88ARFar4JNh9xnTHLMKWF0rZJBXlAfNQu/7mIq97V+LBpbUDJSLotd9KLHkxGVsq
ll4MSmRi8+OnRo6aByuTEuuntMch4lA/tlqaTigRIho0DLD0v+XHfUcFyHzCmfSn
T+DG845xfZ8cIQatO3dBS34TeFCakrn96kaommsxN3AKo34XaxGY3LiYIpzO+pIA
IuaUZP4IJaNysSgeZPhM+1F2ILJgVnGNI8oObLWNYoqmv1mLO/oL7jjzduYSMDJ1
gcW6kOQq9gOP20WLxMX4o0rd6V9YaBKZqqWvMsE/1w3W/uiT6W+yIkF/lg2h7Cbh
8XN/9wwfTTAxa0Jqq9iNt601a662Z/v1fUM1VHTNAhwAZCUsKXAkroErKdcv/9DN
nyBHzabk+nYSWPX7J6LZbSLjXI0eHkFjT35+AgEuQ3+PSKOvAOg+NlEpts/atoeN
NiCXku+hYYhkaIdKq/dSztOQvmiT1oXvmPgMMdKeevxvb4yM77wi5WpnrRVspzzQ
lSTvr7bvWwt0AnyYb1Jtp+PYyiktr5jZNaUJJUVe58cHwhLNxM0swPMPaEscFA6V
SQP5W6pz66zn0Fs8UqJwfrEyi3jo3Fglajwtww+xxMM+M0soE6+fIsYpEc4J3cZZ
NdypJXfs1xVGIvwlgHsozEVn2AnhSV/pA2RUFSCUnb9ZpLyePx1HwF8g4x7+JfVp
9H1WoVFpqyhyVtLfnuKUFa0aixRhMH3cZTRtAqlD4AjUtMzoxWvEG9UZKxu6j7Z6
TOAvQCEb/fD03a6AjbA9q+QzW/8MsFrobNnfayg+zVexJutCd4ZYB7ZxzvQLTQA1
hCOut6011w1TgGzlFli7r/7aFdrI+bzwd531cu+UO0A4y5tiqcgMZ9DGRfSHKQ9r
RrHOLt8BJKZzrDgJDAI8nqV+6XUY9OeS/ojnXD7Ynn/FQi9uBWLWpJfmSyhz2UMc
W8vt0z12aw44Yv5K2BMmAHTxcc5V/bbR6LeuuD31fSwB/1PtUfAzqigSX8xOQX9L
+YMM5DejsoH+R4KIuknAh8GH9crxOHGX5BR6Qw4JTBTGAugEoD6wc0R23+PBXIVt
FoAOu4G+n77hGobDJ2XizqTr9fD7sk3om4TM9eXBYG4j6mjyr/gKFrFDofKaoeVH
0iMK5i96iXk30ClX3q2FBJjxX9Bg8Vb0fjDeaxlPofZElIe9Nr4wx9C1tC1AjgGD
1s2atAsbJ2+iVlMaQxIqrmzDqYoSm5PTtz1Aerh1X9nRS4ldhjI+Nfxr2f6+EXtn
Y91sfE80kQgw3UMznpayskwsnoDK4ZZUCGS68309Acb1BzPgBMnr5MTKNY3WCti0
MGt49KvZf9va9TBHVbjx6lDo2ZHAfG1uoRbM68WdIg0OLK+LHVkYSUUnpNks/n66
wcqTEgnEXCOCz8x75ioiswOiAAA4qaNV0SVTN1AIgroMENPO4Z4kVC+NswuVb6Ux
2q0iiTu33HOwuVMw/Z4LxCh9coDpy0zZS72LMWKoSgEh4IAk0gJgIx0+AdtW+iCh
sMgGe2oJ3dcqzDE5rfIKvjErxD0nar9keUSyY/Ofl+Y3wpIBLOkOFShsmlBdu2pq
gC5IO+TLuzJh56UFq6OpyKtx1SqZuPMcpC9oXavCpSKpdGFFYgwjxp5SkC4ydz3K
7K9pok6K+GYxXIudasQ4Hg75kr+RdgwpNTEmS3CWltpNpOmdQXpywg+wmRiojAXL
qEU1Q4yWkRnmDiiBJplRl1lU6/8EUbzmcIIa89uPKQNu1na/2grWSUF5I6CfXbkT
IYe5TPaX0XDFuEXU2XknGI2fVDlRowqgG+2n0Zg3XbQD3BY6uW+eJ3oc8TN7OfsQ
80U9+f3iYZ0pQ/dSBoXNQ53CARjpvf1tna/7lp264AUjT4VI3eC19G/dzO4uhANt
CY4foN3PfQfzggy/NM2gdWMNDTTnqFN45yLB5v1Pw1dJO8Vm6edmbJsWCyTUBB2L
VtwrBpieHMHuBnQBi5Ch3KilLUnW0vtumMEz3cd9o2S+ZoQzh5dxVgDr9IVnBsfD
Tamo/pz2AbAzoSvMCIIZLV8gYMwym05ApCITjETPDO0lO4tE1/feQbzpgpWFBZIw
5MX1pnWWbTgD/GzhzcqhjkxI7cFoliVzAhiCnvUFSnQNkgXud+MzxROMObHl8hlO
Htw7uQN2wFq04lGXD0A5O7AkQTMQAjflJo4yMBxnptUV66ENDeiEHdV8PkSVWhov
VQs3821mmb1dqFO18eKtdAHZoBs5z44Hz6Mu5v0f8bGZYDZPAa+h+b9Qiw2g5gWY
kUDSiWqZKFXGBdP2X8hIdnFTDkIiz3UEg/GxnTTaoHV6793NlpGG6sVEu4HQYLvi
3bhv3edXF/nxMK2EaCW1KE899jdsDY+oxgauZjakuxN3T5FabpTTyUe9yQM42YTP
TdFNlUY+FX+Zis2CvdJ3BEgz7tmkq6Zw/8MUWwgx0ZF69fc5gkfu60qmU+qAsTxc
+6prDWdfqtaTrnBDCVHyuNc6IpV0vZhbFHRzatB+sGXHCpuiU6MlRHeIybevE1ot
fVnR5R7ghvjD7HnHk/EOVjZzXbo5KXVgis2I8Z71pB+DkNmARScdYvoY/CSmhqOO
BNrLmHZ++eIBB0jSL+mFa8do1fHzCY3Ru5KhFcr8mp1h/Xe1PygI+W1FUc8kvPrw
cbL6XvxwTfyn62LtjffHtkS+a4omhHKPEdNqot2SsGolTQw7pbNkmYYRjoOHPStr
TafLuxnb+UYEjLQOapvKFZXgPoUsPbKd8fFESSYbbTXGXEnU7uACv12IZ5sfLhC4
bsAQJlCOHm/eDdRzwW9kU8msLfPBcPo8MHruG/2M0EvZXSniSgSfa5S8dLBfluhx
G8M4m5z31PKhLq9C2cHianYEUkRTUalRlEJYsm9jlgJVK3CxyngStG2+kCh8XcyC
/KlNzIjJKvRxmgCCMCOlNfdkbmwtolHHKVdAnPHByOB36oXRw9jqlsTSlALErlJG
So3sX8dI713QMAL84OxX+hwgFYyFhg1TLwXDWChoYW1Muy5Sv/sB0URRFrei4Bdi
0oUvxjxdj/euxmNiKHB94zRrL8c5Ns40pdiuNs8J80WrfTOZhAFP16/VTrfaD1Np
BNly4mnoB8pfH6EIqDCWLZ1HoplG7rnkaEi8/HCWXcHE1WxcDqf/sDEMje2Egd5t
Gi67ar3rpSceooCDAAQ0uHf/BSF3/if2xou43lKgCX+gVrS7EAFtr+zXm+Kp4iff
A3xpUTtOt2tIQ4ds7bxx56IeIOjwXYq2ID0yh12wMi/ZeGXOz4h8btVz1h4HQ/Np
qFItd6948ky5ntnrPv4wXJ3LDK5PZP9+qtHVLpevQEay/8MynpTptVoJQPGnHDgd
cWaGUQiwAOGYGrzHVWufDkK/8Ok4XrbZulS69ZJFM+pxfO3QLwD0lKDVfoGzLIq8
RkLLE+5kc0m+4EZcHxKbzfKqyXE3ojzIMT74VgZGdo/vNKrcIf16tNsb99RUNBxE
MSwgQA+xS+sbjYwCx9tiTHFPi6vDm7I/0Byn3bgkSHgLcUxJ/A0kycKx0TisRdel
iH2QWqGgF+M81WZJnxRVDHjk0LOH4aOGTDEMcgx8wVQJSrBgHrrwes+ZXcLzRkML
5x97VUlw4IoZxJniV0w5zweoUV1X665KGKFfl6PlP7dwV2xMQKecO1t4MsebR+jn
Rd9/nG2eVTVbiQtS9332V1ioJjLN3eWO0i3yDX8YYO1d+BakcP/p2mTle6XwAgx+
4IzdkrtO9C1U41UG4TykYy/nTBnf07zg/XSjzuE7FoMOL1YVf2Uwp6+e5H1N/ej+
8mIw0xm5vFyXI3+y1GGW7tDp9fgk0QIewIIGbiMAhqVLQSgj3rU27sRtM5dQJQw3
fNeydIeHWMv89qoNLwWiKTQMDpbc5K/50yh3Eibxx2v9a+tDB4mepmQ9J5VCfngg
xLnYB9v0I72EAoSivnykqkruBiXvTqUpzTrOEkd2cJ2Snyv1YciW4kTjcw299UvA
obtv1lb0RWwMfMfurwAQSzkRXzcUyBnbH8G59WckGXXoEO7jqO/eGNJ1DGK/4Sfd
tr9Si8Lsyru/J9lV4kC8ccvVQh37ucIK8U1JIBHWj7MECDB7/7sYpP5PyAa01hse
+6aP+pAS7P0v1XTSk+GeGaQusFnnraQWKYRIiWOXxPhfoG2Ha2n5fGj597ZSAttR
TxJep1EiW9Dl7TTboZdTkrNcudxfNmljcLFxauTgsKCAjT9XBx3/T1v9ktL6G+ar
bHOu1fvfKfM+iXFBqg+lUSAjNFJIYNHPue5HJqhkCyBhAh3twLGGq8nDHToVOZ1p
tv8qnpdtcL8RiDYfUAuMwmW/CVkpKm7KKpqSiOwMvfLpQOEDuL1fm4sCzlCAktep
GSREMlTn3AvJOMjlzgX+AUqnWf8SoOKULVGsLupPkv60PhxcFaN59Fm1nDtcD5xa
1OCCWIU2qghJpgUGFDRKYYv0+4ZZ/RgbUqtZYb5xKgcpZjO4A/omXbZezowgsqau
xMU1RCBz3GC7h8sgGh6gVus7Sp9BOZNdYWSnhvmIQey8QQMtzVrHaUrMXlEkxJEB
146o1Tx+yRXO7J+997TGy9Z3PLhe1kZJTnSVEjATJLO+nGQdt5e4mn1ZzzPbaoCo
iqEYqiM8LwD6pPPw+hczWD06OZT0T+ua/fA5s2Rmp9nNCz5jWK3wBoMRemN1p88q
i2UnJNZUWs9IGIBKkLgYMBgY/CodGA5qcP4JRDI/iQZnKjegkKDBsU2y/FtpS6pO
PkN+z6e2IuXjAtgsKbgjxpExvNL6wbF07ax2/ubujoV7cpP3MCaXyD7nPAj/gk3b
zEA97KTSN+SaNqEJ/QI3DHq1R7OxI672vMh3N9qSooRqPetcz3Nqtrzolt78boVk
8ZfU225FBp/Yq2RgWGsC+XXJDmC+XrGEUPeLCruBFcoSmpjnAqdsbR41N/6zU9Se
G/fQTpeEAl0PF7v4v92pjDwznGH6nVgPkLqEj3Kki1F8yqfhfMVWWL0yXCU7/u4j
Bgsqla8qJm2LZgKqMHt6Wvlsop3G9mv9NTlICdAAK7e4+r30npQuWfCTgawtiOzp
juUQTbv+Tw5FWF+GsOMOp4+hsOpAQMxscbGxFIrhljlmCc+wTYR29wjcd2SXVGRi
+/K0qYTUDPymXpT8J/EFR07nnHOKMaaZfMl4SlOKlp2Jwuypf2X6uilf94ca8I/M
XAOrhLZ8OOxcxubGSbZ5t5VypFIX2bLa4AEg0vczHpcEwOspnTFko+UhJuuDEv37
mEymYi3mC3yLOf1gu2NZS+ZtE9CCrqBU9MPq+DZdQWoW/26tqEAX14nELcl19yQZ
Feeldxe+PA22cQ/flZ0dtGBrj5BibWCBgpYWyJL4eJfoN3cIn0S1rwT4MmklmzmB
JKOeKs8R2OV3UqD20oyPlz7H8Vlnmu6WJUdWWbnhiCKHHp2H8//C4lr2H/QdFMty
S6E+k9Jvhx+jDwAeBHYVe0b+mkyOgeqAoPZ1LT+WT/Nn6BACWL+D5LAGNq98ow4y
uC58MGdeDYO4DK+XF7NoamAJyuSLRGRKGHlhdl47qVNMf9e7Lng5ows7FJNSCF/K
liFqqKJbBrgcWtadrfMxrc/MmNszDezFrwOWnLJ/k4OyUjrjYPsxWr8oogFxbXvE
TsUe+fWQAH4OMz2T8v94xRi/jKdjaZF4RtYJNtiRclszDDk6Jizrl9JWahOLcuE6
ZzxvfNnm7BSqPJ7AMiLBSoxiZeAHQcz9oinCGkCrYrhTTfOTOe6VK0wtS1P/CJNN
Lk7w/1y912q6sueSRDDUxSwWdFXavXmH11lh/SQkilh46uCVtgO/ZG/HlQS5RkGf
Khk8I6hOkuGixCzA4q+6Aztag/SIgFp8mOJ3cIkUEMDoxrJs9hsv0kLGI+R3jlVz
n2C1OnQLCJuH9ivgj1bj1Znf7f645SEtRW4cyerpUudh941UKQAPh+AmE+pWWpvP
K8YNJiTddRTa+8uoYIEUY2EibfsOqZC82jPO8IzEhPPE8itb/tXyYq2J7Bhft/B4
+bwjyKgu9AOO8/kKpKCBJQKHyGh/PP7BKvj3/8s/5fhG+EqKyK0q+w09CvOQ+6qm
jgdTXHXyvfpum0eoBbGBZrsDSeI8XwqNlGv/pZru9OE13d6xaZ5EbPhcSbA2B3O1
f27TwwQS6fzkjgRZTK8C7R+uYA/8DgW2hxsAQsPBr9SkM2FjxahQPqNcrEYaG3XA
81LGfcaWQk0NBqXpZTE4w81vGLwW+C36Fyik1k8uiHfjjQo++30KiTyOJHG0eIXC
YXHFrChTHIdN0xhaTrsUpH2hN77zGRVQNLMifjWHQfjbA15L/5rn7M2tjPhrAjC7
K8LhQqqy50x85jQmUFtIp4SCj9xDe/eFuc0AHxd7K/Ih3KJH04sx+9u866N8m+fL
lvSWIjJA0Bq6Hic55plUEv9tERFNg3tD93qLxfXQHAFmlRF3yRdZIIR/272WyY+0
HiBFuD9L9lamZk16iTHQZ74PXYdpkOInKv//5slGVRElCzJY9mOaN6bMf1A/S4My
knQtgK6weYYzjO4qOwkk7XQcdoPZwLctcwHGA+ogaVcOyHmpPWWUjcomuind7ADc
g+CDWLv1MpVM+IoTXMXC/DKXyZXYoFLPECMWtCdv8sD2Znfz5ITe/24YsLoVUNYI
70R0RjNuP04wNE+Wl0mM70YKjl3IKIt1T4JK3eZKb18rZDNdDsDARAEB2pRTEhiX
8HGdmEaHNdGSGXigiBlU0DhA+CLlbPT8NRxw9iJXfgveY2HkPj9ro7usamsNN4JQ
n2ULcwRaYWumH7RAX9tNATVlviRgnMxMjpUY7+FmvRmsVMboB3zDz7c9bEwMMqY+
HNEAYmvCgyIsVfWpFe4xDM/nNwkBbRn5JXU/sDxof4FIsdw+V1V52Q0ka+UFzNgy
agnTR5wpF4iGH6f+MUZ9LwarTr06seFH4NohLdmmSNbhJh7SAljTBPGUd3apuql0
j66Uqas0wawc9t01r7k6R5g851Xjr4HwDMjV8FLRISx9IBkBYrTOGd8gBMQhoYy/
+UVCcx2WCHvKyfHO3yVUDxAX1KJzx1WNFQ/pURDeKdduF7QtnzZtnKkDy8TuS5im
2KqHmHLt+0cwX0KqsQIiQmiUrdJCd6eWspEnHQaY4jy0lX1p08cGdXTF28h86y7B
KDhEZi96jE8aBXRq9clDfcGUwNy3n9/Jz3GN+nrFzYdObSpIOZXYOJjHPYW+PPTO
3ALGu2CgGdD21mBWhCNWCDD1/PpmwmyslrDm33iRVxpUSYLlk7FJV+Ggt5IuTF/a
daDDGzDqQAj8zk9TV8PbzZOwgoFU711A3LxY8Z9pYk5pAS/HEyMCtzXPHTTNb/3F
DwH733NWNlxPOb7Plkj5QwIH5OPglYNAcyjtOGlgL8TDPNKVHu6dfCi+0ga44IHt
SSRIA293L4voj87aNWm7BfOtMgde/fkHn/Zifx/kFWaiv5eySDPQV52LsTLWKJWo
1jjd1c4Y09YWPXenPEL1U9OgaQ7kYPa5b0fNqsAmC/zlZXowwLGyLAj2Poe95dRm
9u7Mp/ZiGii7eVCTtYUOfflsRltHeD4izIVYO6hgts5deXebLn56DSaMYjMfB024
I+6YUSnr8mTiZnSoreQLC3NPvWF9wCIXktdrHo+pu9gLUAQJ6kJbeXX6PG+EzFzZ
vlA8Kzj81Fdc/vCTFg0Z8ixPeMtUHrrz7XbD50i60aIe+aoS9pU/PH/2xAnKFTQ2
zG6b2O/E1RqwNcDRkiYp5Y5txfShBlHmBGAOb+ZmJ9ZTSswr5x0Bx0DDy+zV3BAB
p0oGj+pqNxEXjqhae4MuUhsx1OLgfsajWgxQP6eAGv4Uoi/2ugiBXhtlIRzU+UL9
C3eYoc9WJ/Rag/0pO6egWZDX9zk0DXb3SdfXQbcgKgFgTxkjCGScZxYgnePCLi8M
1BPOMuzf65iKt6O59IUbFxbXb7tTBvPhuRK1eJUrkzBDrf21uPWrHBbTauujyPcp
xUGhM83GjkP/r9aCDx1lXHEUEWFMr4uZSB7eRASko7utLlZ6W6mqlOUYYQdsUAN1
ofyC6mu8xu5TPjwj4vhrIQHlpN/vOkJj4PZIlcawHK2T8c1BxbdYkgJ7PdsX+KKJ
ymQe3MtDPG6oAcJxHBUgnT/72TcQMksqKmDOF1g+bNI/xFNVql+nNyOmfMEdFgVu
VmV/4DSNHCnX973/+FmK7Roa/DONoRP3rB7uUd3wnRLHa/2m9ts2OWSzVQAgrCjv
e3ofenXbF8+Bfg11yvd59YEJkDmzZuIBGYezs4+BrQN03CSbNqAyhHWem2t+7p1Y
8HvEpp/3VOo18ywJiZRNtk+WWCMwBOOdon/nhQQ25mmNopz9psy2rHpc1/dF9tZD
T0DJBySqVYEwxXrWM7irjPmDiqA/YPVxN/v/pzTMRSMUWYdIQxSigbzOhBqiVRv+
kGADNbPgcUeCA1i2iM/88i8FBwP3TyxP4CwB+4eEgu9iQns99orpx4DNgbXVR+kX
s4m2oqeiFzSBmk7IZ5G9qo2i9/Silg5dtTqFETGY4wv6UvVo4ufAgXfXz2qbgA1t
wr8R8I93UpNsKg3WcBN7uLihC1fY8a1r16fe68sEHV7eJr21yrCnRr8bERzrJF4C
wrh9cEKQRuKt9O3tOTyy9TsqF19xH1H54vtgxEslJ0BsJSZDiBT1dGUOjqTVkh3T
9J7rCcpBugPE/pN1Jca4a2uOdkPuPGyHbMF52mZWCyA+jjkhZM7Y/zm5YEBBamJ7
7PKbjaPu0BKqvEhO50QiIFKLKV9bNGpUtWWMJl/+iWJd5AkBU94d1NmGLbvbvWX/
Yl58SotUO4EGGDFeHkj7QhuTB88hxcJGSEKho5jRLqs93W8NrxPNULprLlM8PUHF
TORs8Ze+Z00SYZbDCfQqogO4GUy+khVZRMLI+mATCfY/syFkGLRlKoOe17cQD3gN
6OmOSgNBVXmlCvdyF2YYac8qT6JAvbcuO22N+ECLi9Ci01UmZMlsVeVCzdsF4pLp
0bqFb2KW/kPNhLl5BJmBPFFhAn1uu/l+l/+EZ4z3XGEx2/pyoqGWWY/h8LiM2Cru
2NUjfYQ/YoCghxg3siCXWv5kXMgBFn8odnQlJNr5QpeLmI2TdRZnm5GwawxWmv2a
11jhWTchj9X1LK6V8f8CI9nVVCQHujYi1zyZX+hObSHRriAGb7fwipQa2lLYpDDv
2+c9uIqbDPBQInch3vUnhR/ZvSlLPyg/YVfzPNOnGPo2J7uAxUMjAYddyZiBa3k0
A5BCJmGcuOwv6PX1v1f9rbkdrrF9AXFz55ry1PHyFbO3O56G7/Cx5gz90gO50PX4
u8CO92Bx2K+hzOl2Zg+BCgRFB8JZZILubud39OYa1TdVsdlWEsj+fcrhid8J6utx
MjgvM3gsCE45xqblavn9Pm1hLaDt/dS4HF32wNiY1kOAbWUrvVLkCvjiKe5ZiYrx
BcgCdRWe81BgZAgGwfQVIKA0NE/cmUf2wfYR9/KsWqnjIuTSp1cO6I4+B6Pxaxsq
2Urt+FP/X3XXjioq8SE4/9dERIVKUUUyaGNOGCYSxMIVEce2mk5Q5HlQQrAfoI3l
dMFaCKP/Rxr+eyELNxFHt6mNP4UpBwFxfTRrNIJ5pVrxStUsDYFakUysaamKgNOa
Ya1o+elZjQHZEh7y2aV/yZtzD4E5+M6pIhw2JCy7W/3IA4S/ejFnmZAe17aH/ieL
gAfE5d0jOwhHu+BpRLzxepF+xPHpMGxvLV1nGlg1spjDLEebaxx+eZJbxeF9H8Mv
NWrDFwEFOdvyGVP5VfTR2wwz6IZo+oSWEbfLMIv2Vw1Nc3FsSHbkc1CGDnW8hc85
LiJs/9th730q13PqVcL8C2zkJeAMS6QAjVSXbFOZWnFPcG/w+zPvcWXD33rysFzw
ffBsoTVWkRvC0/DcvYjyCgfGt6Jjo7Qemer2E6h+OLxNgVIBA8IsQmonNivdiseq
tFYsIKh7BplUF9fYAcehVEYDFA/HfMwGn8ghwHeSk5EeD1GkpNepukiTAGxj1cFf
2ZxffpyosMIiXvmEnFIVzFpAwR8HiI9KkNdJTKeQKHefO60pSR+xC0pFMj+aO2tH
RQaxdCObLWqHFdIkGP7GIoK0Xz+O6mgw5dwZjL4PmsHhbyb9g3kWzO5pgaAAfGHB
2I2yDfUipIvaUSHvuNWy1g==
`pragma protect end_protected
