��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H������N݆��Ȗ�����}������XQ�ǔȀ�wu1eH��F �O���6���5ig�a%���5�Ќ6\�f����^ŶG\{���6��5	��p��S}��jO�@m]�;�ˬzgv��4�i"�d-Ψ�C��2�g�˰i����xW�2���g�~�E<�?Up��%����
���'඼h�{��3�%r:���r�A�KL��^U4sUf�])���PBf����ˋ�n���h��OWT�LT�9�K�X�U�k��j�&�����]��=����������|�)�
�3Cu�	q��me�� �ȝ�C�BcTg��,,�%
�#�6Nu��[;K-F�n&2�����}�{UA%,z U�>���~��7r�zDJ��$a�[z����-�~�O���~,`N?��7r�:{�&���ݲ�Az�WSsk�۸�I�Bh��m�d�~�y�H[U��n���s����@�Ĥ��OJ������jҵ�u;�<Y��7�� !��_�֠z�hm�����o���z�3��,�[��xD��~�{F+؄ؤ��߲6�ocW�?�>��,����̿저_p���*i
�A5D0��a�TbdG&�1܎�>���q5h-�s ��7	e�^Y�Sl�?&R�� B���ơ�M9���)�s0�E�Q��^{��K�!55`����-yx�����
�9�HbcQ����W��f�I^�թc Uq&Q�h�~!�l�o<}]6i��N�"@�P{۾�4*�G�1�
d"�^�7!�ʎc� p����,i[�e�sBH�*�I9�_�p O��&^3�܍[s��ZGj9�V/\��jVRo7QI4�����DO�h~��ǳŰ1��A�w�}�:��2�8gw}'�u��3��L1zmOi��
����Ԋ�<��!��4Ymh����^��]�`i|we���|GAŞW�=��������R��g�֏�Z��L/?�GK>�ZǦ
�
"R��?$	RLX����K�H '\�㕚���pnP%9T{r@�d��*�!A�1�2�p/f`yHr��Ww&��&)���g�JD���c�r���o�eE��[��6ܰZ��(N�=����f3��a��O�U�SBX"8S��lU�
m����mD���:��'R�/�h���>��7��J�W�s1��#X��Ǎ�����kr6
�X�U5�W��vS�D�.��z3/�@}�^ы����0���S/g RV�Q���	�u�ܭ������L[H�\^������>B��(4�n��5ʢsX��Y��!L�I��n��/� W6���(�YHn��f �L���O}h+1i@r�!i�Q��>�$�Էv�>K��y�GO�b���������
���k�]>[����)yH2I��3��Tm��\�w��l<�;������:���-��bxJ��R���Ef� 
�V���]��#�62�4�2�k}s����g���jG^��M�f���$�X�ƘM̙��� ?�����ҠuD^&�[	��M|>~�闊�b�4��cR��4H@YxT��D���O���T�ǭ��r��r��K�~�?��6�<k������#�u��w�Y�ڴ�����쏠nu ^k�V���R/�p��
�`�_E�}�c��ǫ�?æ��Erc�n ؿеj��Sfwt��͋[��4�9G�`;~M��ta�1~���]r)�$(H�.9H�_�^����,�9����X��t��눻1d/�����Kx]8��I��}2���Z����,��("S3輭̓�P�a��PV(�%����h��E�³{��y�K�XņS"71[�ft��)�B��������?�v��r?S�y�r�>߃��@�ޥ��D\s߅K�'�c�j���11�$�2(�G`�3�}`e�|���5 ��B�pO�PDˣ��	�@�F��c����mp)&t���-��cV��D�^��88ܠ|�՘1�P�S���]}�Y�$�V )�(�TC:���2�BD�}1�mB�gI}GzdOC�g3,A ��}��ᐤ�c@�e�QY�;�"�0v�	+)z$�x���'c�ޠ7#�w�I�C�:t�]s�s6�c��m?f'�	�"
�������S;����E��zOeh]����!E�G�1�G޸�M<�y��,"N�܉nM$N������I\3���ƀ�[`�W�m���!da�#�6���u��	8�"R��g5.�:�����<�����{߀���էQ�H��z|^�7B�-����7hRB>���&�/U��Ur���;|�2�"0�So�����	PZ�����)/R��x	��L\���.��.���VV�^'��c��]Q/=�R�"y�;5��z�Ǳ��F�~u��߯�%v�Z�[u�J����M�����?��1XV1�����w>V�Vy�-D9Ω�iz���&P��ox�߅2���'�����yoF<�}Щ�P[�TN3ƅ^���~!��� ��}�u��e�M��FH⃎��P��Nt^�u$Q����"�2����g�