��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X.�84PT6�3V��ou��Uެ�Μ��)*�2���y��7�k��Ȗ����_�H�U����51�� 3��
��	�l��\]���=y�GQ�Ɠ!��!p��՘H�\�%V�\��OZHx�5��.us�H�Щ�\���Y�o�kf�e/3q��q<,Q�K���k��n�vƿ�@�ۘ�3p&�Za�x�|El��9+bBS �|�aT~�v�D�"�]7fF�A:��wG
�(u��3�HEDL��$�{ r}A��z�8ԗ��-)M�;�;.�zv�E�c(��|��5^��&��\%�H:ڹ�'!X�QY�E��.��$�#��|����� m�I{��<Q�xlq\$4\b��K�8����'��щ�o1N�ro��Dpc�K�V��'�2,�d�+m��?(��|9��N�*~�04�|���>Dy_VT�>_�Ff����ހ%�#ev���7���^�j 5�J����#��X-�9�d��4ր��I/d�cΜ����t��M�ztm��*��}-��C[P����'Xf׿�y�8�1�"`�#�3�\��N�۸Ӓ����.�Xw??ƺ��ʠܤ�p�L0u�cl�=�_��,A�$�`��t`�
�jpY����g�+eC#��̛���-��r�)A��)��aB�b#�5��!̱����l��h��g<�	pl��W.���\�5������q�3���(�It3<%���%s����'�>jU`�A��~�!t�=�z���]���1_��&O�l���i�E�Q�bL0�-�Q�HGE�*Q}��d]{ ���&ǻ�~��8[���ðu��8?:�&yᢨ��Q��!�d�1+;����>��GF.LMk�'�Vw� e����4�����:�\�g�UD��%<de��XFҝ1Omj�4#[�&a�(������'U�v(Q*F�w�.�H�8M���*1�����@�0{�=ax�EP1����4�T���>�3Nn
dr��k���ɠX㰈ˣA>�ܽϵ����}���喠��F��5��\ 	�dj�<�g;��2Ǽ��	o* @�����O(8@��Ĵ�P��<C�|*������MF��^w��
���1�Q�ūe����}yH��ҳ���	r����Ţ	�?��%9]p~8-w|1^\F��`L��;��>��Sl eo)ֽu�}~]�{g
��V��m���՗JbQ���U��Q�Jr�%��4Rs�"��(F�MJ�B;�
@�[�*h���W���X���S�kA]�+m�n��A�Ha.|�F��"[�����(u��K�G�ZVw�!�/ٓ�����=�������!�%��	01uC�b��:m��3^!���^����F�9�l�"���L��+(br)��Oڏ
ٖ�zB��W���Q��cGcG��2���{��;UH������^2�F��l1��ҴDR��}����>w���\��X��0�r+{� B��^f}P!�L�k{V0#���;�t��g��M�A�4�����?e`Q3��'��6�\������_�,@}���1�Q��G��*�c�&�w�T� �F��t^{���9���*ŷ8X�d�`�Ѩd��`~2������;��l�Xٞb�c�ٚ�'1�H����t]�ԋ'�z�ok�{sE��#�ﬆ�X`�>�l;/�ə��h����kJ�}:�/ڸV��+j�լ�Q+O.�|ՆX���8p4��U�K+��F@���Qe���t�M �wo�l!�����~b�@��)�s��F�P_d�9�f�Ã��9��i\�b�ldW8�wxA�ra�kb�5��J��i1�{=G��g���lu�~��ujҖ�>IK�n��2y�
`֢�g��ҥ�Z�	Q<���	7���h?~!�-��0lg`��u�dP�@�W&�@SVR!�#�&�P�#I}Se��\�$���ê��#�����7�yM����L4$���⪊W% �Tq5&��8nx(v�^_ᠺ������T�:�e�R3d��*ؠ*.Nu��	�	�X�>�=�t�.V<)WP/�غ��~W.y�ޟ4�D�.�� *�d,��o��m�:�J��]5<G�獱ry�<43��ﮙK�N�x���G��k`�n��&&I(왵m�%��Z�	u�(�B�d�_M4f$/}��ǸU���,i{���^!�8�K+�Cg����%��4	~i,�@ܲ�|��������h��3��o:�ጔ�g��y(�td �Г� ��:(!x��M�	�J ���s&j�.�V��+U%��?������$� K���ǝ�t�0U���ߟ����@2e;vA�Tt�q����<�1��1��a���,�!'T-�'h�ρs��)������ȼ�^�N����q�����/L��\Ե�z0��a��-�wY��D�^�%�N��2L���3��D�:8[GC�� �Y�t�$PQ�V"BHw�u�ھ�4&[���D.�oӾ�/�]��㦿��ޗ >�_��÷�x6�D���0[ǩ�ΐ������a�9[��N�O�X�L��J�h[Z�����U|�\�9lǆooɫ�c"�||ה3����IP�LiF�zE�ٵd�
KGfS������H���'�g�`c��d�M�3_� u���ۙ�Z,��XE$���o�5�`g��q�->�Q�*qA���,���sJtc%|���ozI�Me�� �EzO8�ߩD��ర6�5�s℘��M$�xM��#]�t�q��^��e+�q2B\I8���`m�Np�q���e���/�Q��xok��v��E~�����D�p���_Y�1e� �CuD��R�Mӈ$E��:�_h��$�#jl��h+v'C%F�S����Z���ORS!k	`���_�W��f�:����u�6�4M��m+���zN�)1��AY�~3�RWB��o�E��3,2�'b���p0znyr���[� �T֟8̡�W����Ͽ>����0��?�;��8�J�&lk�)�d�*qʅߋ��E�˴�T��4�z����o�OS���1��<����̫P�
�(�Bq��*�%<����J:*P����ܠ3@nS~�I�d�»%{6� �2�d��wx}�~h�c�p�l�U����S�kٛٻt�E��<�^��P��/���|8T���yih<ow��w ���c�/F[�S���"�x`�����}�c�����#�������8�w �r�9eE	i��φ�����"��(/9��J�h����b�]$&�7#-̬m�H��`�3��s�!VĴ<^��BS;�E�ic'�L����<�<%Ku��U���P�[��M{*g���X��<0�
���!\i�.��q��*v|���C��^�S�s�  �)�A�@� �&�l�洝�ל�j��c�;>"��@w!h�P��Mc��GӔ�-�7�nz"R_ �t�[��wS���d�@W�b��C
s��e[�!��|��7�@��8UYp�M�\h�|��}m7�?&���SWa�c��0V��TȺ�Gh u��\��P�/7���0�H�
[���-�/8S��<=�ч<�_���u���vÿ�������[B�<�&��ϟH���|��6�h=tG "gz+i��s m�� ]xY:��~$5�2�tģ�w᷆=M^�`(=���ղ�6Q�~{h�מ3��e��a�����K��?K"�<�"�>�e*�b%��gh2)Ү���l�v$S
_����@0+��D_e�����Vޜ��%ױ�S�k��} ��M��.���/d/��5���R�#+Նt����
8�p9����-�'g��qƭ!V3���S��Ÿ"���,Nc�\�^��HB�R�*�)�X���G�B���'E��D�r?P΂�)��Z?Lг6����_�"�n�0�^!Aw$7{�$�8�+{��t����k�f]����C ]�݊G]�F��0޴(hU�:����Qֺ��q˨��qр�͠���YO��j9ɇ��G�l��l�\�ʡ~\c����}��b8���/�!�(U����In�d&��<�"��T���P�&0;�#�Xԗ9��Ӫ��E������	Z��VV?ϓ����<�0�!���"A\���Ch��I2^XT��x������VDy+[�d�2��P�窻i���d��5^:�Um*�Р}A�5��;�.�C���|"�� ú�ţd>�ڀ��"��H����s�)�m��X1a���Vܮ3�䵉�ȷ���ڼ���"�w��*�U�ş�x�ɡ+�)hº�WD�E��6���xv�{igi���G�)┩��y�,��TU���N�h�ZiǟI�Z���ٔ��-`6�m{�/�� xd���z i	9t��|�[�^Ơ@e�@�&'ڄ������!��D(Ň>Nƀ�+ �����zf�qk >�ʤ�b���
3[��g)��u�3:�'e�P��U޹���Ǜ�jy�F~	*)��������l"�tF�z		�.F#�,6��F+�>��f�7���*���=�1N�Cެ�O����x�S��Ow���E�E-T��M�(�)8�Xǌ�h���� ���Q`��Zu�-sW�͹����]����L/�������n�>k�9`��{�ZEm�X!iE	�7����� 1�حV����F6fY���]���k�!������?H$�L���"%�,[t�D��!�b���e�EmU�GB�b���%��[G{T���Aȧ��,cPbfm7��m���\�B��? 	�g��Q6�?d�)���^Ѣ����䨈�d���=kC'x��G#~�n&�k1�K��2��4E��Ȑ��bs�b1�oj�q���%+�{9o v7U�q�K#�*qw�q��#ޞS��ye��,|��K��S�n�2c$�	U>ҥ�L�J�+Î���SK�ޘ=`%M�� h�"-J�����E��]=�I�/.���������4���K���9Pzd�4�	�wޮ��#�]����������3u
*�PD��Ju�+7_��Z �c��p�B���ahL��å焹!O��d��>�wtgܣ ��M+h(�����w"�G&?�q���Lf����?�Q[�Bo���,��:�c/#<7��f����&�����}w�n��0>=X�-����K�z���RD*~1[�_w]��D����,���Ь�=şN��.�� ���؝L�H�%��S��*��A���/5����f�ď�^AXh��)gz�BVw�ڲ^�s����{X��Ǟ���.k����ʻh&M��PZD�Y���vX���

c�5ڮ���T`��1�\>C�(���U����7ck�Q�X��9��{��;��>� a&��f�'��M��.��͍R�5�J#l���Y��*���·�=�����JH#��Ӫ�q/��hX�:r�iS��@'�p�B�~��l�]���S-=�W�k��`͟񨞌x�)0�,�U?f^�K@�wJo�r��r|��%���a��|�fxDN��1��Q{����?;}�o+_�4�����L�j�T8��{M��v�c�Y!���o�L\
|죳��7� l!��"�z��T���4�V
c����]OxT�8�Sa�F�<��x�r#r��v�o�nEM��w�"Oe�it�Se��\���dq�8e^8]��[�B�Aa��������y�m$�-y5�ċ��9z>em5�q����~~	�è��hl� FԷ�
u;~E®����8�|{9��c�ٿu +^��ә�ѺC� H�o�5b��(�7jr�AXW�:�e*"w&�}��?"S�����%��
�d�>$���锎-f�����Z(��玌~�X��\�G#��O����U�,� i�s�1A}2\�I� �Y>e�v�Xe��o����,q+��E��Ts�K�4��}�+�}J>}7H��T7'��l��5	'j��y�Uic�P͇��I<��G���{y���C��*�K{���aʉ1������-dL���x�	�q~�[AG� �$Ьq4�n4��qhvTmaoh�F�z?*?���V��y,�.���q*�<�3�i�Q��lp��k�6��Ҿ�l%Eځ�x͊|! ���<�M닅@q�F���?�yM>lFn��&�*gIj&|��K>�k���O$�D�ڦXK�װV3f�O�?�٧���θ�፯���d:FCo�Wl���Z7-��	��E��
�Q0�`�*�9���2e
f���p���e�>�N��$�����!]��n�%1�s`�i��b��QK=vD��u���F51v:M�"��4�},T����Q$Px_g#mvk?���5�(�Yh���;�u�AY�T�~�L�q���zߏxzUA��En���A���&$9ƾ�5ҕ���NP���8ΜY��¥+q1� �ƃ�P�ʽ��~ܫŋr���҉-�~N�w�1|p�E�\��F���^�j}[�\��蘹ű`y�w����=�ڣͭE��D#V��lD�י �;�d����(@uA�Y"*FD:��}�قXg侭ͷ#BG.�T����k�����ǳ����]�(�ӕ�4��P��B��s��x,_O!����j��>�Ȳ�%��^���d���~��0�"����|6}#r+jq����Ue��p�2w�{v{�j1Yǵ���� .�A����ě_pքo���&D}�T��!�T�I9�O��W�ɯ�1|y�VD�L?��ڱ���J�H<��Qn����t�l��tU"�Vl`�!�xjXԨ��j&���]mr)1�8�-���>�����/���#4Q*d�)مj�p��3?x�zm�b`�����.R{��̋�Ӳ*���:�)�*�R�8�@��8~ޗ8K��_γ�����2�a1����i�q�.�Rԭg��`�α��ꥊ��E��:�c�x'�UH=~�������X�;ln�1tC>b춪����0�]��1;�;\�i�P�:��'�Bt߭K� �%�p�ng�F�Q6�)�+y���4�n�5���K~��[��3��~%<�5�����2�gx�7;����91�J0| =�*m���#=I�zZ��۪�����?�^H=����˟��ܯ��^��J���D$��ʗ��_��<�!�O���ԉ�m2�7ʿ��=�x��a���HUB9�,"2.',�����>�hM�:�G$�f\��u<=���҃X��j��)gL��XZ4��U���9���ݞ�&�|��4�����1�W팅�����7���D�O���$�?	0}�_e��:M�:w�RT�qú�!|�:��cRL� 'G�5<Qh>IQ7�T�wtfD�?E�EV�ZЉ<�����jO�Y\��`��h�.ǛuX*[�Dy�z���.k)EA��[����^��Փl�	��"g��ʱz�z��hP�YLݪ�R��hGz��l��T�i��5Z�+��{G����;�򋟟fژ�@�6D���?܏��B�ٞ�4R��J�Bm�詞�څ���� ���[ޅ@h�K�u
U�e?<T! ��g6(�ܩ�1wQhf˷:@j�}Z?K/�����a��}����?7�i۱K˺i�z��!y6��j���kP;���ԉ��O�	#�A=��,O��ObÂ�+���?�~9WT��:��r�!Ĕ������$Ys�5�X�gK���A���?�r<x}���;	������*m����4�i����=�&f>�9^�G4*����2���0�#;�2�k����Ա�\r���D_umv��"����s�W_~K5|)�a�1��/.rK�F�#�W"R��C�G,�bɤ�o��gu\07L�ZQ>�k������FW��N�S�	�������F�>!�Fs�v�2:�5�i���ŗ�g��록���M mCU��qv^�=���r�	E�����?mv�[��|d0>���K �'��9I:��z`�|�I�
���3�^��'�Yi�S�݂�ץQ$eZ�`�UJ�x�A��ʽ���������-h�Kc?��R�C�y]K�V���s���JV+��FiVh	_��!��j���d�wP�@X��%	������"33-k�ۓ�S��-��ɯ@�ZS���� ɒ���9+L�VB[���;=��v���ˠ`:��&N��P �7a��Nv�Jn���Zѡͷ䃥��xɖ����m1�F�q�s�IQ�"��`�����ɟ��mب���\��L'��z5�ў=a�9������y5D+��{��&R\��hf�Ţ��r`�v��D��*gx�G�� �����*6!k'�ꅠ3_��Nm+9yDV>B�w���qS~�J°¾/��Al�d��%��d������t|�uo�H�Y�GC�0����X
r�8[���uW�s�J0�<������Iy��PI�;��"8�8��z�8e�悑��kGvK���e�P��U~I�(����݂�ţ�sڨy����K:YJ/>����r7���b�5.be���%�Ԗ?,5�$��t�=��~���^����q0��Kw�����gE�2��;�tF�x�4�-ϑ�+����}����>�տ��%��[�{SY��?9���Xb3�=eƖNe;󘣧$:�����Q���6���e�C7=Oˈ��� ���)��<��犩���k�H���
��XE�rd��(���>���Q��|�՞�|,Ac��*9�=Ґ���,V��C0�"�%��K1������v�~��KS�-�w�׸G�A��|'��	���c>/~f�f��b,��5�+'�~[��(p�<y�R�T��IԲ8���p��3��*��~�'=&�,/��_)ų�ZkX;�(���V��C��l)�\| k�<7��H��;��WK��YR�ͲY�e�U��y��Ф��wd;峜��j���P�g~V�q�Úe^�2eׅ���A����\���*1�O��Q��q����MDVj|�]��uz�z�?��9�q�b�)e������-P<�sI�&KL9�뇉]rO�`_|��ޔO�%��%�� ]�� �J�Z�4h^UX��xR}���w=A�����#I^�O�ү%ע��O�޷{�ôZ>K!�ᨑ7b���X�_�S�\����-I��A 2Ӝ7e�~豓F+d�S��3O�Z�Ќ�V�������)a��O+E|"�iа��B�8��j��[�!�������NBL��>|����h{������o=�-iА��,�I��x��N�T� թ��~�s3FŞ��<,��������ճ ण�V=Ȩ��c�'s����:Hi�p����c>�ް����W�p8�,'�76���~�	��pĨ	M�>�z�������F�=��.�q.d���A�L����q.�C����v�z<�2�o�Z�S��Η�l�z�i�lO�T���6dy�0Q��^ �9G��fY�듓%�Z�>Q�K2�h3�G1�V���3Y0�}�p+?�1-p��x�����W�'о��+��]v��9�i�������.��u�`��n���WL�D�I��#�=kx�ۏ���C1}3#:�c2ߡ���_Jב�a�=��M��3&P�2���>��۲Km�J �Ss]E�]N�z6�w���u}jz���R��:K�Ѻ{^���
�ɥ`�:���� XP����.U�a�w�y�P��G�Az�{��CB�ð�f:%/���	D��H�Y��l�1d�a�z�ޑ�=�q���ݑ{N\��OtMa8��+��o��(e�V����s�?xYp�匚�A#�_�b�?$HؕÁ�v��0L�Pbp�}p�`sb����~.��{�K�㑚e�j}��p�pf�����l��$�USi,����Gl�*�D��z ��N��̯ؿ�#`Q	%���6��^��*p��(=��]�NUT�R��[$ӹ/�3����'��=`� S��̩Ѻ�ƺ�]O���Q�Ϥ�pW��9����T3
��ދ�a��;i���!C�����{GX��Ώˑg�,���Ԅe�fl�*�\���3�R����ݾ�Wn~P��?�]C�J��(�m�u���U�js����m�	�-��̱ܸ���X��1�����[�W�� ��L�׫p�P+6;K�Hq���H8��jҧgXG4����\.2�p���_Iշd� % ��$���W_�~ײ�J2@/H[��r���&0����E`t�M�B�i�j����v�~��!��ؓ �`\ߔct���:��4¯�R�������K+�����P��w-:*��xԏk��\��('z��E;߂�OC���8��4��Q1A���$�2�]��װd�S�sgj�����^Sp�n�|}V���I7O�h�5d6S����6m0�����Jn
���$X�C߾�t�5��Z��$�ؕ�,ǃ��9Ǳ��sn��������%��V�h=�S�L]�����5�Q�G�$�瑼W�!Q"���&���f�Y�O������zJO�����i1��L�g��~�٦�o7Mf2�T�m�L*�!3H(���F��Ђe���e��k$c!m�Ї��������OZ�}�	�"��Z}+�(��i	3nEC�E��2��#�h��]ή��%���-�;dZ%�
��|�7"nācS��=���MIl������ �2F+��U�lH�%��Px�N��,�<�gn�����m$H"�u��uZeO�t`�4w�]ɐ�X�i����Rj*�eƊ);�&��\��CR��5�t|�ʹw��p���B�?&+�.u8Yε�Ὲ��&%=M�C/���+��<Vc�	G{:��N߹x�sɫ!�L��0n)pt�{���.�D*+�P��B)��p�;ߞ;#i|]ú��\ch�L�09�0��U]:vY�ô��w�R�9���gR�Nф"�Cp���]#�Ry�ra���K+�8�����I!��S������mЦ1�:.�� 7~�U�����{�v�;�x�7�\	_&��|�� ǣ���&��A�I!��>�&���T��.e�韈�i�\��.H�4��k�I�������n֌�{�b�����f�w�ʏ�:�N��~��M�h<�؟dE��ԁ~�z�9>�����|�q�<J��h�<�J�����T�7���l��c����"#���[��!-�*�B�ʘ�_l|P�b7�]�"��r��#����0]�&s�l��0J���.�(��$�a#�9O����b�4(��*
=��K�0��IѢ8�޻o��QȀ�ei7�����m���9���0�ƠI��Գ�1CKN&��\�Cyk]���t�.��
�ݨ�Y����R	��ڔ������;�P�}���;� �jĈr���
�J#x�C������C�%+�r�m-��K����Z���Ȝ�{�u�@�[�t~/S�_6=L�75�\˰;�n�~�,s���u�R�)q�:�O��QF�)xB��Y!��YZ�?~�������H^�f�g���ww�Xǝ��T{^���@a���ͦ}e3�K�H������K��O6�c)pX�Q��G=����U���� ii�2Q"7�{�4Jg�nܞ68���0 �Me�B�F�=����i�;l��(1=b��s%���(๫U��j?��F�����̔p&�*R-��	��+��F��
mXs���]ρ���Q�2���9������EhC�8҇�����N� ��A��Oq�nI�Y6�h�@�Zf:�3���DC��"��-���]�q�]P�s�@���'\����,� �
����,�� ��7w���'��H\�aѧ��Y衡���BfV�bQ$�A-�r���R�H!�����(�A{RB�:�3�V�%���O�o��mR��I�=���9f�#�q� ��Yl{z�Sv(Dպ%�l.��?��N�ʄ)
�rr�F�~�Fh�	���[P1 S�'�̐����0�R��e�Z�lی7q3�<H��o���<]!eϪ�8aˏq�cXmU>C�g��E?y����E$�t�"q_<�c?(�E����6�Q2������?����R������m��G~���{��(.K����ϩ�~¥@�Z{Dr�)3�E��@r?MQ�InW�-�W�1M��j�p)^�ׄ?[ۧ,ɱ�ƄY�4�Q���W��Mǣ�/��VanZ�5;�
�}�ϱ�H�'C������!�?~�[���\0�}稨�������g �#/Y�M�I���ŧSn��KR�k;�R#�g;;XJC/p�b.��߸�a	;&�����aE�#�*�sX�p�ڿa��RV���`�r��D���������cyP�����(7� ��X��o�x���aF�5�T�SN���y�U����=;KR�Wя0;����=rx�8���sL��M�ǖD�=���4�GL�$��L�{T���>���/�/D���u����0�h`�ѕg���0�B�%�iV�t/�)=&��U�=�O����/���+C@?�|#O��A0�-�l҅G��#�w(�Prl ��K?h�5-��8�����C����1�2gM���]y3��Y��UP3���zُ�t����E��^ڕ��h𐾝M��S�0T�f��Q���Q_��D[@�Rc��"��Skp	�$��Pi��JY���E���^ Α�N	(��dH��[�-ԟBqnl�杨.8�;g]�[俣��.�����d�5���v{������+��)��R�@)֦Y�8��7$�m�9���"p}b<L%��3H�¼pƎđS���MՖ�L�[�чYZ�p�5�P?7'��F�S��\�����i�q�~���ţ���ǇsRGi=���e���^�Ht�?<a����'K���r���a	���_�]F�)��
b��}b�_4��X�z��d��d��r�fI�xz������iÛ2�@�œ�NFa9�t�f�f�5��%k�c� u?4E���1��I��/�l��*a�Q���r���n�)�F��"���ߺ9FTR��3>a��9�5����:O��5I�))l{�&���.0�rFKz쵰�O�8�i8Z"������o��;|�!��^��3��������3V�݆����Q�3h�h�uQH.�dWoc�����U�cޝ�.]��|�-s�������� ���Q�*5��Q݇���r�|*�&�����Q: �ؔ����N��Ғe+F�ņ\��d"A�6�ȕ�2�ԟӀM1��AW�"�)τ�戕:!�w��?ć�xw�
D��S�Y�!�i�.Zsx�T78�Mx,@�ƃ��%�?�̙\.�r�W_�fY2@[��c�gxڡ��[��$5G�6~d�r�4ց���·FC2�y����E8o`=�e����L�$��3Dy�?6�'�H��j��~�%j�Rޡe��}K��S�����j��A���g�21i�C��r�{ji��|��F�a<�TP矡�&/�F9�����H�h�,s	i�,�*�&o1��@�����e �upj@�A����ā�Tnu�F��d��XjW\ɞW���D� 3�Q13䳱UZ�(�Z�G)��MW���&Q�|(8w¨3i�*��ɶ�f�ZvP��k���6�>�5�	�&�����$E)~j�=-+��M�S9*/�dP�N�x�	UA���1�Ā:��jJ+jb��ڋ��Y@�f�AW��WؙsG�@L��}b������O��zP�_��}��{����+�w�Y?3�І�;u4|�g� �T%'J���O�t쨴�p�Y������3���{��e�W<�cfӺ�qA�6��Qf��!�Q�'Ϝ��Fk����dM�@�s܍2��o��2׍�Hk�X4D�����Wa̽�J�!��FDv��շQy��5�?y7"<�2�I��/$�l6�&c�_�U���c<�9�}�8Y����"΂�6#��g�[i�U����{�6�NC adjMW�:)a5���-�V�0�D�A'3�]�	�ےH����x;�"�3�3��N�/�����2�"���4Nz�C���N���)[��G�8�o����$����4��w8�u�� ���O�4�ܭ
�6������\}Z�~f�U��j?[���UV�� 	G���K7����0����Vu�E��z�nת�gx��E��J�E}3��6��z)S7J�W`�N�>MV�h�^�����u�[X]�ν=�.�t�^���~��09L���Xͅoq�=v��!$��ˌ���:�+�H��V�ޕ����L��_
>z� >���Gwu�02�n
���?f�C@k[�����B��{�D�H�5ڢ^�w��B�?�k�0wg{��i��7�����@�C��j�/�ŮVjK�x�}���A��piJ�M�Q)�0:�B��YA��|'/+��G�aÓ�∏u\P���3�z��V�H�����:Qd�����p1�*����jv1[=��1�I����JT�����V��x;X�����+4p��1-,~��e��{�T�9k/�xke��Vo�AJ���$ �e���11|q�zO�Yf�|���-&�L��	�%)���B�a�h��%?bSz������m¦���|�'�'��R&�W̗�,��X2�.4�� &@��γ�]�Zy\��6,�zeh��\� �R��HEc#7EjJ�O�f�
�-��p2��k��.D�.���R��iP~-�#4uL����"#�/!0ӑ@,�=|C8PN�{�S�Ү�}U�Z��0Ψ/���`��ZX�W3ѭk������3jS���(D��0��}J�n�P��j�F3067��DE���n]I�ȏ�����]�x-��k���޴�98N�IKhԆ���[X��W���z�Ӗ�XG]�d�����/ӈ4X?v����M�~����1�Re���@ `�kyDG�̠\@�o#�BX�M�= �Z��2f�q.������	I�jĞ8��b(^U��8F��v�$�i�o��7�1Ê�S����^��.��(�Hg��s���5��]ȶ:r�a��8���4�����Ʒ��e����	h���r@ *�g���%�a7���{p_́�K���?�
.S!��Ϫ�0��e�6�¿��=a���e���z,�5�uc��+�~
���������G��}�����E�	�h<j��9�%��+1ý�'ԧw`>~�Iaq�*K�=	�;/�J����_8<�h�y��Y݈ r��J���ʟ��R�5)ͭMqlBյ�஧�*�JA#j?�#�@q�L��j!�B�9[!`R�Q��Ywki�`c�;pH�@h��O���S��G�^ $\���Oۛk��L��4�qI�^�S&���tAa�Y��I��D��������٘���Q5��A�k�umԼ$�lF��'rI���6*��j{�Ҵ�۷����w-���L�'��ŗ0���H�b'4�&�%Y��s{ھ+	6-;���B�a���s*h~Q4Q+:���_f6�cxp�yQ^(.:V�L<�u�̎=���2��嚫 ��C���)��-��j�P���<y�[�aZŎ�f��*�Yjr,��gQ� �`��0 n� P��![��K0h�37״$T��:!�� ����E<|���( ޶9��!&��s�wCi�(�D��ǪrX{�����i�_��#]k��Q�{-	a,�醹�'nΑ��w��ջ3F���Ou���@n]4��B���)!�о��Rw^F\�|1-�l���/z@�{����-����fk��63V�κ����X�	�3�h�?���C�Ր������
m����o�GU�B���`�4:���1?c��d����U^vv`=���%@�3ZD��]E?��O�a&W�	M���J���Ph�KT���`�E}�7��?k I*dI5�Qҹ����J"b.�y7��S�s�=?p����_���P��3�D�0��A�DAgBH�-)'k������t��"[͆#�$k�h�n%�b|��e��SQ�z��R��_I���	L�ݦ���O�"��Q+H�c�(#���)~��Ǜx�<[�ܠ�N�A�h�d����������p�,Q�<�ذ�����o�BcՄ�n@���2�ڟ/�nH^���hw(��>�z[��G;�>��ނZS�Ah���p�a7^�z����k��M��nruS1i�xCl�	")o79*	�
e�^Ws0B�`{t�������=xb4 щk��>Z2`���d�����e�duu��g]^�:f{�+\�O|1�����0���u2��`�LI9LN�E��H�f���L^����g��A��*܄+,�u$2�|A�#A~�/hei�ox�44�FO�^��;���k$�u�JV8wB� j�RJ#��|�_�g�=j�b��P���^����.!�$`���.S�Y���+6A�h]>Uu��b&�0�a��Qdq`�?�7Z�&��U'Κ�'o�7�J[)x0��# !�i��^�����C,G`�߿jwt�L1��5T0�G4����s��O}��f�G|V=�߅u���,�R��YG��7y��R���~3+^6�����6�����sK���G(�}t�߽I��14Ŏ�U��qt�>@>=T���#�s�0U�P':�q'(XX�H�<�������.�Hd�Q���	賥l�F.�L2�2��Ӓ䲔<�gVfꝁ�4w!`�����+W��#{�����:+J�Uu�S5ǉ�4�h^8��A����r"Г�G��%�����=@��L���A�p���FS7_4ޞI_����_-{�́��x6�� "�DF��`w�Y(yoQ�Pג�����|1�K�BǨ��DyaK1r�FzUb�gC<��qx���k�k���a�f��QFD�ˑ���P*۴�n/q�h^�D�߇�R"��/�O�kP��jQ�w�OME���hZy��[�9�M:�!���"��p7<3�%�����~��T�,ٔ5j�� ����KK^7�Jb6;
�9+��6\���������t����w���L���i�V%S�Y&0��Q��:�3=$v�XVp8�:G8���j;>Y�!�<��eVū�`�LʶT��7�ɢ|���{��N:zm�«% Hgr�5�VQ������� :H���"e">�Q�#�QuE@ ���_;R�x��O�կu |��I�S��/�S<�F��K���_���)��;����Ȱ�M����������z�>�>�g�&A>��kڥ�E6Ѭa���d]ݓ��Ф�������_X�N��=^��DW�>ج���Q]_��ZNض@�Y�
"��#���7�yJ�'�����Ǌ\7à�L��������_?콽�)�0�O�;�;Is�r�%F&ϙⶽ��R�.W�"�Jfl�~��t��N]jBd���E���!U��|��.��'�d�ݓ?4]�0�(��;�A9�+D�?��� E��T��:����Q>��Y<z����ȹ�����Hɝg�eñ������me�L�� Mm=������j��	���]�U�*l��WIGk+�bDV���Az���D��JH%	�Z�D���]�Kyp��*n�xRg1o^$#Ǹ��WY���nj����S-�M}���l�^�?�i_��CQ�e��'!�Qk�Jo�;�}�k���-����[�,���z����)L5ǝ��f�`&�v��l�~M�m�U�e�W�`��I��5[�v�'����������X�fA�m�s�Ev�kM2Fi<��I��[�z&ƶD��Y\���h؀�7M�Ȥ��x
o[ox��ӓi��b.�Uޮs*e wLjo�QJ��69=���t|a�GbQ}�h��A�f�3/h6F`��v�ׄ�Jol�I�loY!p��� ~�B��t�{24�Kz�W��(�M%����"��rqi��TyS�p�\�*�KLvW�)����B/�J6c�a���Q��5�!�L,�R"ٌ�p=�M�zn{d,אUr ���R��ymaj�z��fۻ��3��ܨ���'�g�?�D��^Z	@Lӱ2�B[4X��[���-+ӻB\���5��*)xV��HY^�RǶ�k��&�8�E��k�4֍��ӫU���~�
Q��$c6�oK{�k[���yh ��
�|��A�sb�!˞g���"iF����H}�,Ca�ۘ��I�e�6����t�'"����N�Ł��gcy��ߧ9"s��:�8TJ�;pY�TZ�"}H�������p��_� �@����
�(�.�J*f��`���7L���r��];��e����hd�g¹]`�>k��N��j'�<�B��E�w�J+���Y}G�W>�s����d��K�k����J�ʇ��'��xOw9L'�nSWȥ�l�Q��ef&��T�3ӟ�F�N�H�|D7�{-��BC��0n'�:rz�U(�.���ɱ�I+9Y���c#\Z�v_XgC����$RȖG+\���U�a	�45V{��Ekj �2[c۱�X�dl����'��"CDr�#���*��L��eVow��B���^Ԕ�bT��L��׭��	��l����N|�"S�V��^��P}�3�KjB0��M�o~�;�Vg�3�rM��� 6#<��m�t�����U�`�C�2hAj��ʛ����{u��k�����?���P<���{f�*<M/Z�l����eO�B��%�6��9�@�N�
��d*���#�ˇO|fl�����|
?(�d0.C�k�'���S�>���o��?�!Jze:�I�)��e)A���JH�M�����t��Y?����!_�iM]םPڍ�]jIC��h�*����_0�ͨ�,fL�Z����^:w��c���T5돚�l�? I��z���b<ѪU��fMq�)��%l	��U�y�6���� l�  �rJ�9���󺴱&��	�>[f��I!Y9k��k�M���!�4b(-��o����$���yu4�!*9��-!��G�,�D��R��m�@k=��\�C� �ڨ�3��`�3H�I�W����L�Ԓ?��G��n"��B�s���m�H�����aH}3#5���3�l\'�!Q�/xPo��??e�S����� �4�Iǒ��1Q�x+�^�w16AWݒ
���J��ќV%R��d���η��Q ��g�]B�h8���H��)�����|�Tv��as#j痫�x���c���b�p&�%�q��(a�����	�`��(Ɵ&ѹ�S<y�c
g�@��.��S?��]�C@sH?o�5�6�����@�����]MN���/{>ڲ����,@]!'���UB��^�ߠ+�H
��0�70ٝ��[���`�+9����Z����/O]Ws����;�?,����j�X�ԤHn5N�β� ��jF.��L�����w_��:V��;�[��������w;�^E��*�[ {�	��lG�Vvf&ǩ��w2Kz^!%�5C)�Z���:�hJ980Mn?���B���_F��I��'Xw���R
P��?2)�/!'/����ޥ��/9�k�tGҤ<�Y&���	�3�n����.h�Zī}v�����8�G$3/N3�]˰!ҥ�^�Gnڳz�L�+���6q�UC�lE��-�"j��f(�'��')���e<(-8.:��������-#:PÌ��6��2��@[�C�;��^ �P�ӓ�����F�fŶI�m_8[v��xx$^H,����1��j���7�u{�Y͆��0�T�I��v�ܔ�x�؍7ы�^�L�l�؊�^Ak�߻�Фt�y�ow���Z���4��+p&�S�,�c �7�B����Q:��ҭŶ1�|1�H�U��H��"a������{T�P�N��
(.�,��I��A�%�����*��s���b�>ȲY��$��r�m��ّ�Y�H�2�.l���)�X�9A�D�n�y�Q"�����g����*�S;�n�Q�E��=&ai��%�U����)[�04���؍�C䯒��޹y����Vh_�ԧ�j�	��F'�,U�α�My���V��Ԏ�!��W�q�Io�\�?Rɸ^�>�9���]J,�GqfW�c�tsU�FKj�T&Kg�-6s��M�2��)��~�|���O\X���� /��FVq��s�7�� �1߿5l���ςZ�1f�^��G+��X�N�N��י���f�0�����ܡ�<J�X9, �f��3oG�0.��j�G�_D�RD��gP;��Kӭx��r��I!�wzC���q胖.��a���> ��	�V��}�㴚||թ���~�юYPG�ݮ����2dzn'& �5�\P� ��&L�8��F��g
AU��(%Q���Jb���8y��Y��� � ���NP�+� a
���9%K��4+�m�q�C�!	i6�B��Y�0��ɱBy7��(�ٸf������1}L�57�d��,7�F�,�$�]�0�B������f�n�&q˰3ڐ��\M��B9N�m�*Ȯ�L�� S�_op���j�\��x�[��q��P��6��ƭR�H��B���"�8Įߴ$p�ֻ2���/�*���>Ŷe���~����wb3Dq����3{=[�$�E@�&����Q���D�[U��cl�hW��a��������q�(�˓>����%�E�~�gO��B(�Nu�o=T/��K���+>�/�6nI��޼�m05���*��C�(�R���[�����ٸGd����_S�No2�r�F���t���*Y���瘟��R`"��fVVU�nڮ�9V=k�!n��)�!O��S�+�ic�O�*W���5غ�m��|H�O����[�<+��r�]�Ii����E���1�/�0�q��[e[Kw{���W�U3վ�?�~�s�1��E��,7#4GH����C	=z��p�1��.#3Af��N�HK�~���~\�?o��Z���L�i�Bt�k���C�8�'oo�u��M� �Q̊���Nx���s�>��0K�5��3�����Ha����&��/����QX8z}��VRb�WLET�� |i�U�[z���%��a��DD��؛�0�W�k?0�	g{�#A�Kf�8eH��SJ6�'�GA����K�]��%$�X�mgR��ͻk�x��ji[O�h*�@s�����ۓ<�g(f2Z�Hᤧ��ڤ�Ai��\u:Q2�:7�8�j���?�ҒVu�'�[��E�� ��H�^�S����l�,R]56��̾� ��T���߷���r�d�c�B���d/��R�nGM�b�/�z���?�Ʈ�k�r\�/;��,ϖJ$��[}����{�j��*�|:�fK��K���C�8�":8��r�ڂ��Q�L��M�8�����X[SC�>�z�J��H&P��z�_�~�3��e��K�u�^6��R:Ժ� s�8�GQG��27�X3�p�h �f�j�v�����Te$>�(Hh�x[����g�-��������8n@�H	��jdZ�:�v]�̩v��"�i�L<~N)���ˇ�𬠶tՓth���PDc:^�y��GG���t:#�9������m;��x���2�{�lh"�/Tk�u[�Z1q�0�������ڎ�A�+��������Uv���`������FוL$Ig*|�T���B>,5ujN|�'e�Yx�����㹂�Hwq�����hI6�[�p�O^[;Ȓ)c�����c��E9��lM�O��`�c��J��d�n#��+/��4��(���o�Y�2�ĠD���<LP 4����z����U�y��FXA;
�c	>�I��-��->�~������:�"����o�R5�*d*��g��f�_�=D��S�z(�{Ӹ��ޥ�4��isd*ӧ�S���=�m�� VǠ�e�ɗ�-�c����2���k �}��<�?�|�|���w�`MJ_4XW�˂*G�r�ngT�14]�H�W�=�U,������'�n�/��L"��.�����s�����5��~�\)�P���!��x#�;�m!�5��Y��RFTls	���6��½^9"R�wI�-���h@��Җ! M���I���O<8�w����*�I��-�6>`G?�c��D`�<w�VK��  &p��6��̍v(����'����al���Y�J�$�]���f�]Mc_9�D�F/~��� o�E,n���Z���ܔwΜ�1�1��iol������wd+@*��GJ�B�y��Q�4���g1�O��� ��Ŝ��/vV)~�C�r���(�犙���2�C�It�O�z�����og*�$��gR�9�������Mڰ�qn�2���07��v�{>�G����s`�3?���%f�D��S�����p`"�4��sY���Z����0�!
���Ԉ��3q��ۗ�1Sj�ڑ���q��B1�w��o���(h��>��N�[I���S��<?JDZVN��H��z�C�f�F�B=������[!�T�I�@8tGr_��f�|����[�Z�m�yԬ���X��Y��gC