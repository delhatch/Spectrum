-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZqK+cv6W66a7LG9GELWCyH1wGHUekjn6xhvUj5gEnW1vlolaTLhUsTwpMCxlcnfWYOkK/tGY9iC0
M2soawBNra0pWLbaO3extwp4skN08YbtokL1X4nitvEZJqR4QMxHlqm1eBidAK3qoEhEjdS3/e3Z
CcjcVr1GXo8IUmga3axPVMxsBvIEGcclhDpTke066cgzXdaBIQPYzma7evqu8JsQnjvmeIbjefS8
bNiVArAmAKjnybm42B70RJ9fP814XiIROUuSBo+h2g0dK7t9HtyPjMJ71raEXzMX+qoi87tGBWvY
KaIJNfcxYPanXoZ74pfU4Zf8QEwkzdlQx4vP7Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
N9kx8lV8r5NyDvsBWbIg3Np01MhgkY/+DUulE3KzdnpSzgVvc1YVNLq1V0LTyzbLKBMvUWTEk+uI
67OHJWeIn5IsvdYDwy6bQC8uCg0gmxEraV2eiT6QhS8hpPtNYV1EdVGD3A0pxG8IvB/nqYin+LAh
m5qh4Z6oWyWOSh59DF9UYIXVjGDl8DXBD/yGCrPYml5wgdLnxeNSmzU7I/0b6K6K14vcp0zrGhmM
roEMj9XXgsH38+qJNJYpHETTiQBa6IrSVFe9cYjVz6n6L1KlPKaKtSUhvYze/lG7C3jpUWjnebYu
Nm8MmtBdB2+EgWqOG1eSurUhl8stA6z68cUHRBGxJaz6GDuqVrLUhUBd/lSzjE9/OdbCCjM6dIqY
/d0yg28nG65ujtvlZO11bYyTO1t4Ka97ea6Xk6ZwA7GWG1a04aRzjUhCXWh9XP3nLqjltcEBIh4T
N83FlD1Wq7dIdXAwLHV6iGWpQ3qmT2UrCt0fXsbGffxNv4kL0ac2PKDWylrcNTiEv0BnrNdo0S/V
ZV8yZJjJ+PPzSuNUaLSapoLkvAqKBVVsAd+WvcTg1gzjUhs5xcyLt+0nypIgjRLSmmOY+T/t5bNB
MHuJ4uLTFdI4NbR+l32jWwOrYOsojzwZUUZQfIPlEn5WPUdNpNIQK+L5G1LjPqC0w0r3yQFb2/DW
aqOhmKQ254ZQxrahqLBdscWPidimsj/rlcsPoGVps8KIqnO5/I8PjZfa+XzpnksHtJ9QSKsK/ymj
qeV+N9NR9hm7mv+aQQ+a35CqfFPo752LQNRAsuN5lkFy2ikmzxF8GL6/oWgXj3phCGny/wxXt6ZZ
1TlnkMBhlmjxizgurLreNaFNe0BXvde+Bu/ld9NgZNWeCJ9Qe/oZRDMYiIln9DjwoF/aSdFyNlzL
5b305I/oGXNYQfdOE2mFmPj6KgYYytWw8Pv0eyJWtXQxAaIsD9sLgFMjYSYQpkMxg0qfev3sjdcz
3dvXxo64hDhAXkJ5iL8Eb3c6aPWo5z3nXVa0R7i+N76h9ZwmmdFnNlVxjgvMgzfGkEcOSkhHhz4o
T15TWDYRTSYrdkPsWYan432WB8C6sWqmLT5cDS4/tnWUYHFrXtGO69dnlPw1fo8fzbsoPp5wDDpU
BGQAjTapL1uI7NJBhOiufUIn0FfFUij8H/aJ9ldJN44sKwFNHkc5UkQAYTAns3Rf8MKD5Rs375f2
/oOqA/Uo3FP5cGIYxvpFy6MYX2ZxRqLVABYeXd1aFOSHBCtEBvJCpQfAZfdRKO6tGnWEsiyxAefZ
kC5cCZM4A5D6HrvVrQNI+/4Pap570N8wjtRb55jFVd1BFAUCeudDPmEli+y8Hu4musUlNPnv1Fun
/HmEt0piWcBZw23tpDP2b7Iyb1az+W9xd5abk28n9u426Zn3gCDPqtscBLGqg4Q9NrdxGRAATF4O
mjtdf6dCrJqXYJSXLSL/+NMM5gQI5fHTXag/g3tLPKUq6FFXod5OVUPhn90oSXUEx9S17ZjH7UlA
So2xOIkoI4ePB6llp56YPKA3hPQ7J19/Wbszuwrh1ja/TOqhTA6mP7wxIfEMDUYEtHj40RcJb2k8
ZPmJYof0ADcmMS8EaYr4d/jdCPGrkqdq8hAvo5jbn5/iMv7t/dusnXY41bRIa3JSpfRJ+3NrJjTa
jvcbvLFayCpCeG2jP9bfpt7JMPT8cV1d+xsC+HxWPR+EE+SC93gJkts6o0tLF1Oskbhd+4GZ7Twl
O3V1frWsvz8cDvWGzDRwgbvsY/y+EvhRq7COYegblUbybzTJ6Yg72Yvdsj/+MYXly7vl/IYTnFuL
QQgrybzT/Jm5Crhh2ZFMybgQlunH2ezitRdU5aWKxn9Iy1TMytZPPJ88ommRe8tHgq03gI85Hivl
wwxlfiNxnZcxNnoCAp4DujN6hkfAyQEKqcUDz/5pcsvUP5qj3rv/CR4SrXw7cpzcOFFUfLuBPaex
N7SRKGNN1BAwRHe53hfE4djzBzqXvcsqtk5x3lVqhJ53DEaPmEkXOQsX6T1UyY67bmtVDkv5o+yc
e/6vgHKt7wS9wV78ARnClhS6iGAc/uKv5NTaaUICHefdTWBgLpOZVoeaSt9TvaepV5t2NdVcfvA1
s/9+f2BxYbJh1q0eRg7fD9exTBRPnzTY4I/8fVt2SAcuaFcuoprcXS4+BkygN2avzDANO6qynERv
1y/gd5rfX0vFwBbBKJGXsvN7VoARabHTGIKL9v1KHiXPymnixIodZxFqR8NbJYFab/iS94noPRy6
Fom64+mUgUrTyI5TsbVFOydP43WuQtuuaAwJpqVOMAJWPw1gFlVQd5bMFto4uz6rv1TYE/Z8ACke
xRyce5Ubgbh1foEweeen36qcGPEdIFpCJgDSK7elV2xb8WSWuviXypjox34DjX1QGE2b3M3/w5be
9Krnm+WZbRpT766ynwU9dwWUoyQmjq+IYQ+etxBcWHEGr23xy40aZheB1+vX98Wj8/z5OzA1IJ/P
np8pTrL4TRD+2Laf+ZOsNaU2Ts54YBwDGFynbST1ep2wPCK4hF8nsdNynxLM+guWZmz8Z7drMlmw
Sn/alxOQXrWToac4QKl1HX0fHFl/3enlY+zfv4nxYBB0O3MmwyCkgXSp4TFR3eGYEieXYIoeXNwH
ViFv0pr/hD8KduZ2kLLOKEWAtIfbyBVxZPlDd5u3WgGRaYFHYWGfLQpBa6QI2wgkmBBDQQ5qG7WQ
KTN2nj5iIVYwKgu7oTAp3SqNGR51DrfJDZlZ4BJ3spaRs91QiKkeUP5AqN2YfYt/2wn5bew2+BSY
O7rLTvXDplqsfWxtXoiMQPOcU/G2IJdZYObfPPQBPbcea2QGt4CZzqzSL9Rmn5PpkFiiSrswBrBb
NCDQY3pZuyqgqnJyiqa3JlgUo8sXHcBpZfZQBPiNGxgfk4lUGE5SRd3pW/jI3/e/1K/2TMTITpbR
SB7W20NYat0MaH9uwjAAJLMUw7aF8RHl4zOrhXz7o8WKu7lM1RKtup+4RGBrR2Nalxek6R+//qQ3
LUro8HQZNgXVOHjR4V8URnhThat23YUmHkFAFaP0wPlBC3JF0WATbyl5dJoDFSjI/59baPYBTs2i
1OLgZXneMG73TjKsg5IqHv3cXvKDPf9D30NuV/czzquhODE3T02u9tfPOESs3w+2OImFGhqY+hKR
QbSlL/TAtXjHQFF6+w9W4CrUXy/VIVbon4Xulcv5WO3H672y9UFQtndQRnR5Rx8n8oRVAqQfYF53
Mu5YjzCh6bRDegBNmJb3O+YnPGlFzLh+eon36aBpCV7EaCI2Pb9q6tGUATSE6K9/rS8OBvcoI4xS
QqjehigK2fdW9R7/QmAmp15EfTTk8YQLDwtjqnwXfSuqyzfa6eByM0A9lTls2L9mLaW+6o41kv2b
SGq19degaQpoMHuUNY9R1M8mq6gtIte6loFW1doft/9O4uEpliN1al+TsNPyFev75+uDXL4hjeKk
mMRGVWl32MWvzPxM7+Wnk+G+ghvy/PQKsKdFZsMp+QnAHCAq2pyVGHPM+nM1Zummay8EOi9UMw9H
HSHTBd8r9KojotZKGw5QREo2GfRT/gk4qPnlG4B/V2vBvjZ3x5eFhW2V7NAeIIGB7SbKVF560j46
OF2If3uDYw71RtIuPjsVbsDvlcX0Q/jPkBqBDDFpaCu6aGvQKHSqCfqmMZP32sTAGY/Wrh3I57C7
tBq+Pw2QhFYArioqLL0pdZCuVFHVbIJvluLFAGawoQ2mB9sL2de2vHH2+qkuirf8DgOdHnGVTEH6
FUkEA6vLLEBOGneqTTpRS98Ro2XhScE8056Rdhl4Cy5QloFKCKhOlBVW9PwdMKq9dVDv87I22ISL
gX8Bl8rSrnldQLM8JfcznKMy9vDoTLIZY0H/zdXoAp9xsCjstpe9fadSR1tQ9+QOxzLVTSqO0d8W
xt1UAkl/8Sy2ntutj1i5hYehdpxWs06ERq8M/DvN6U9/HlvrolSKMwwPkWEFsWLW1EImHDjNqtHb
JwZTfBaWazIfJiNu18sJVqtuC7yv9BeVUzwnhV73bM0eQo/o4TDVCDVoStTjaLddqAt0hZDqcMSS
SFLQ/Tb5nHj6L+Covv30wL9iDioPGe9/NnreTaKjFccQPrPmXLXVUh3IDMUO7CGKVwpL0goB6bx2
1CicFwMKc0FsxGk0qxGMiqq4wpQzS4EQByodA3i8ai03ZIAaoO+K9OkTodw8af2wca5Y8LVLy4YN
QMpoYuyyHPl2LopMJHZHqF5OPPnm5WJhURSqlHn4sU4fLpONEk+Ki97Y5mCimPSzWlyQBceWkRXB
AKwaeEyX0pphZO6hKi8ALda8oCbpAPIAW+46nh5QuRmQbxbElVRCWP78Xm3aNqRGitB+4BtC88ip
i8ta51erE8/3zYzq20wTRInlKlAWBqvQj0KRNSeqlN0uXVWWOYm0dI9NZM2y7Zqxg+D32877n0lU
7RmgLR6mTmAG9EyW8a+d8iZHAJ1mkNe/ybNJpzCb7Txbm9gjZ2YRFstGg29ILrzaWGXEf8DDjAnw
cuamU9yxXN6rJAQl7IZaMztuIdx4HwL6OUV1JSgb3GcduesV1YsVnjcNIr/90KLkniQA4PQcdGvs
qhqNnVmA5/iZiVU+uFFoBIzVbMNAGTH1xkYTW7QdyeMEqOJosyp507XIj+sRlq/D5wWJvrP4XVzD
B7LSRRPMm5ZmXXHA0R5gfUNPonlzs0IVTgY+dKDsF/DCU8WDOmPQyl3zW9qEM4RIXx+ujAMd2oyx
B/hoY6AdXeXobU4LHIfCTs2lWtVM89qKD8fcq71i4rvYHKtlMmUoGJeg0Kq8P16zipUqhx/99JKf
5jomaN4+cZP6u7SQ7uIGN+jX0DBrLDP8Yp6PZ5fCyPHmRRdquaFRJMoKXtIAKGI5l++OqEjBVpUY
sdVYRTwUYvM6aYN4KomuNt4IEQES/RKFZNWLWgShdd9yAnciB4pPvI06kzkXEcVI3KQzduHdXz06
M76x0BrzZvP+vXVVpKofco8+upcEH4uIx/xNKjq5mFpNJmSsyQX2eYPFRnjeKVK7R8iDeSHjNxVj
fmS5u0Q5JEdJK2OjdBnkj47kKfqRdyep+nCU0yGQxzsRHdISqi7KMbOZ+MnL0qfGnwqWu/2mYiDQ
oZsS6sLxHFFR5YgaYudewVRsT/mWA4kjbAcmVW//YehIVBgBq++IZ8T1uPW7xdmmbk0SzUq1PmfE
P/Fl77ZSb6R1UdyGoiWfTk4pMyADuSUbAUH84HM3uCirbJQtSAjlinYffvttDr60UlxfVSElnqWz
6tTPWPtHxzZ77IaHqjUt7DfX2Ml/BdtqUbfXI+kKahS+TXrfaU9I+w5A9IPeSzvBFLgNbC/655w4
GzXyJGQ8iPbgkgu4MnZ3wjsoLfVg/mCqi5Lqwda55PSP0ljMZ4MxjrzaCmdj8Wq0Mv66Phh3veA3
Z6HtFFMsn11q6ZmE1yVj171Dyes/CC2xsBg7s6SvSCNX5LYoYdOv2XIiWP3aRTEtMqSCmBo7CDIW
AUb4FSC0d1KLYRYxo7PS0Z2zT6ezvwTPlKHHTLIbg3wTaIOUCwD3d4mUGzs746qDAnimsSd6LwWM
nA+Ln9zbnYCZE3vBj7S1WM97PIru8WU0nVW5n82L95XaKTmJZJicSyOa0gWzLsfzz5nJGljVpNtf
iaS6FLuq4A1tjFjU/brQT5AZOm+7KRQC7A8UQ6e0GJTqnRhGRPCoJINwC1rEE4ysffvqLG0VasGP
AE0obXxndayMWCxyjuQHM6ql+5HHnEyPShjQC0WHaGnJX0bGYCfEE0gWIj+4AvBiiutX450uI34D
MFHfr/LacS1ajpkB+5MKWWh5YiaJU3Baiy0KkQaTWwQth+kaLe2WxcwZud5aa7JucC1NnimTL91i
bRc8ClA/D3g4g2Pf4b736NFfMbIoVWsf1zYeMWeRebitMyPk7DVlhG/sWsIR88oW0TCRddx/a8mk
1qd/x+riprEtDA5gWuzPbZqqW2ruSvnsPPoCJrKpcO8SARPUs6c1BfWtjSvhwnZLfhbKkrDIKyIY
qpLuuaUSqRfZQHAbgV2p1s4mofso+WI36eJm3eww0UobiPcLBZyT7KXvucCDUUW4YtH8DXKKzfNL
XXSJKWNk9ATIIfFNXi2w+bdkWpAyqhyKiBD5YMqcOIzg4ms32foogpdbiI4Sr3p45A2wTsOEqkVE
52EJgPDes5slmQsHtl/3wpGW/u38GOJD/Y6x8H2MkqG31j4SU2Oi+LzntalWtkFLbgRz1w5Wl8oW
vJzn+Tj77Qoav/rem54KZef3lgbTFZvoqMWozQRnZhdPxJwAfXpXSgwnkWiqXOmGXvXpbmmBDEbV
0OxGHZA1GcCbxjfUajxk8GqfTNJ72I56xU+LZ7AkhF0jxU1yFWV5GVMsN0ilY+X/qZQQPFUzMjTQ
VHOtN8dNij+SPdyVtbhSkuMhA3ngfpr7M/Yu7ZibzdukzO46HWfIU1TbWJcfhKqv7Mdx05alrqEJ
1wDVTzaglP1c7tp610prVBgwX7fQAQ2eWXgWPgtPyreAVRGVqF0gW/YyxlN9wTGbdRXHI2wOfn+O
CVfyErNSeQrYqJNMYOSa/nxbdLRRaXO805GmZK8OxrOTW1Dh1fWPEjSwHjFxeIjWdziUfNc6/7e4
I5IKjW4BGvhf/lHnINHoCUfqaBLXA6dbPlTV4ePRiS/4ym3m/+w8FeA+tOE1CFd0BaVvSCYnjFTF
iG1DHe67Qf4wZWWomiSl09c85LYfvvn5wxkJczfBufG+YKOswjwWSXJgBXlBmV/tWCQaEOq2aBFO
18BUExn7Qa8VKPXCyrMhmEqVFXjgiE6q8aZh148s1LgRLxist/zpfo07pzSevaqEW3LV4heyvT2T
sNRTP7PukXD/ceVnnIMrb+WwcpBfL3DyzewyCM+aSzyTBxbAAIK8kZViOpTNy94Q+DmJlToPz8x5
lhu3etYwLmkEe76icL2IkDm9B6WH55u2gH92NpQTHhW8g1UBHh17K6HCvk3I+en0eCvW0FBy4daa
H983qJebG5Kp0i6h78oYvqciGYO0rM+COnuanJgFpXJMzeaGtQSryKgQDvMmylr8qMO9QqGFHAbJ
/C8wQtAAvtrqLmnqBQMYQ+DKqChh2jMNipwvOa9YesbWdx5zNM7rVCATws7epnEnQPbfwNvtSqP3
d55IpIYvyrU21Hd9Gv540dZDDLiVP3+0A3mOZf1Y8lGjtYFqX4os0FPA1kvUiEUi0TaGJnVGkDhv
PYLAkiSSoQdCJ6Z8K4m92d9TrUWbbhD7C/8xUNqY6Xd0wdvX04IzezFOUibmbz/5LkIIW64/BJR7
J8GhcALFH0jlTglwRmwem1t+LUrRlySgyfwmvBW8NAvY9Bjyqg5kaVWeRFFw8KNVrcLVQdbcY7MJ
h2RP4eGsBUKoy/Jlwjpc149rI3fN/ndR75UC5djHPSXi3OoMPvMRaG3tbwmCqkSfYhc2redHU+ec
fCRDox5Fik0iTXEGMiQZwU7YGY27vv2FGUUgnYbvO1gu8gOcXrpr4NN50DG7kImVoBjMiUhhCXqb
VNKMCTfbzXEX5GTwyd3gCHz3kuf3t8wac4CPzRiyLy/PVh0+5lli5NkBWj6oVQIxnRmJrN2um7Op
I7+AYeM2NNVE5PtXk27lgkPO+FZXmJRX6iGQFrJnOLWaaewaWc2W66vR/OZBiWwM8k6S6tMW6QJu
j9vbBDqwyCSZiFvKucsbQRa64IIe316aLhJTASrDOqCABlI8XESQKunmzbClO30CJT2OdKSkG6he
htsJVhFr5eTKOQ9Jnqdwl10/w8/ZsOlPPglzSriWO2McRm1IymWWcGHBeVNC+HmvilgRUg2nIzAs
hKv/mLPT1UItVAe46XOoCEFzxWRwcIJgaUkK0JxeCurAPyTAaXB6uSaMw6ibSU3x+1z3Jt73NEPx
GSRrmBb/wGsgnVNI2jMNY9xcTTtxC1Ak80KWxfELOWjC+sfM9Dp85ufN0E461+tA+35rut7GDVJR
sMyWCdDQ7fI0+wZF6yBKMs00t+Mg0VahlmGtNibIANJf/GKdE2MXfVdetp+MfZ8tRkhYlzalCEOM
h3hKBzp/p8MJ5eNvP9vVFEtqVmYjep8PImq9YoF+9CeU3t23wDgqtCzPXsYpSGhN3Uy0V0G6akPl
3KiImneItmXJxXM6pzUaxY1Jqka3qepIleSgQHRgvC89zDJ5OmanaJmGEr+YujIQDEoPMhM9FqAP
oPxQ7dKZTNz87tt3Ez7T++EY1Z28mX7fV32vD1y+QBaK2NXivqzkkTJYCOdkH+7p8Zw887xRnurQ
yamfHqdbBXHC687V2BNc/XNYRlPfamSIi/xtAnAoJ6IfCrZnJJutt7bWgGyUCJQTKUiJn+kSXejD
kcKweGVAAqJ3ROyyWwpiNeL6JYbZ85yastKRCwJoWHTu/pBqqFQEpOvU6TlOcJQ3az/x7XoxEkQ6
PBiKZ0GSaZvnCMOUjiDYKrtYZFT0OUhVBItRii9OupvlfnypAdunDPPvyBC4t8qRINb9VWnEsHrb
5alzA9/vjbZvJnykkTiDEhs34K+g5Sx1zsO3RoZ10hSnouVSQE57bAV9UjZnC0tjTuTN2ohgFxbo
x+ekvON1P4aek/sssiaEMbeDdm0ddO2N+bW3GaSxsB1l99ZAnxH5EHtDY1Fe/fAWRH1eGIwmT2Pp
w7TyZHa0z9UUC7CzyaBAdmCIKtQYdSO86lbqQghhTkHlJk6nRu8r3E0YSWDCnfmdkm//xfDt4Huh
Ft/1U5823qkkBAPw1JrRvG7ePmKRZhi67kPOWrpB52IR6vxHCNAGqYtLVAc4UnQW2PZwe/1NxsZd
bvMzFSnigxAj7VjsQtx6zPPpRBbBW1QzfLywArw6PWR7VbHyiWt0TLQ4avtCJuR5PhFsx3udWrVD
MbKi8g++pDB7TSmpU3uynlciJImdkjauXddMtg6VPoGN8URbCB9ih6GDgZ/xFWSnjK20Ewld0TfT
R+EB3OorRxQTTzbBBtVB5Zh5hyaZFy3j0PUgnWdlcp2CKvc33Kd0/jXidPPvfnTgYKrw48x9qlJS
iTbGmf4I6JEfE3LK6ZYhNGYUiBoeiKDuxsOn0UEcNtyt3mWmx0n652I5X9VzR/PJYKAGybg89DlO
bWUT7ZD12UI8syNG+KaWAMCBKaD7YCo979XXFHV23GWZzJahaMgKCy5pcrxVgDh5eZBaeuau/iTQ
HqPUO8tFAEAqc9LXUvwfAnBs+W+b2uG8Jn4yLov6Pkr2lKhnnrHC92iJHX60nnLMSKWUpHb02OXH
LI9ZDTMA0bemG7l6jEk3EC5N64YDg3Ma6GhVjl0GMTSr6Gpg8KJyW/QYSTjkTPvfZSsL0mdQcdoC
TV8QlpQPCPM8AnJQKJL7amfD0x3w+vJuhuC7BZaYW+MwSCuh8FAIKVgU/GpTPgjvu5j1lOdp88Cv
vWM+DlYL9l9g4lxhKgOLAlNknmXZv7wIxPfJqJ9UWMrnVIzJWW3+EZzihl7rWD+/OBl8/xHlgOte
EsbR1A84aUzV1CKSmuPeh2WqMPBXVn8lPrA4MKRpoB1udyJ6bBlMeCmPOGhm23Ii/+awAZTT+JpC
KROGduDAqnyWMfJ0qhygv3SWZmAcKvsqmvdFZ3TGRxgkelAtkhneaMZw1PF4+68DDuidasctplBW
qrrNWcTW1PUVgmh5hH2GbLIepU61YVK13FLWMKNMjhRO6ufoD6V66toc7Gt8JvhTYt1GxNCXHVHo
j8vC5T0iwLTvNGM+lmp/fR3VgfFpaVfwzEMHfQZkAtWw24FCvzhhQx3Ol6kat+1QAus9Wv3iSJyV
A+AoXbMtWpI7KvjVSx0peiHSen5AhHfLBJJC3+9pGfCNawIsjZ7PcjGUGyspKZj7l2LZXP9yYTQ1
EHqslBVKXKNBlMcDebcVp/5edr/Xx4+QWRUwoGMCd9gxKDyNlzyvu2Vh6kMo0BZfLCreYRCWKLZR
lDfjgt86U9qanQstTG5EV8hhcGsNmfGWLTZGX5sCO8x6Mhc2mwG5o6vZGP+iIS0LXX+p8Khq9UYH
PXTip4174lyijivPISqMD8FruhzZFdRWjIZiy+lha9JDeVun+ie9peLSkdMK1eg2HAWcEIxTx3Fm
gqY75YkEx4yyUJ45NQUrUINEhKwPsFVq0cqnmqZnZ+kWjMrnQ9/gDj2UHmUyGCqsf3xJMqzHx6+1
fUsnKmEuOUoSSU70J4BIQgnx5GQ272/XbDNRhN7CzCX6TY/aLLNvraYX3T20w9JXEGSImf8lPtER
68aA7Vvjn2m4bJMpV//kHzkMlkWfPAnqt9ueNFSaraHRJjEC4MdOmEYDQdyVeNQkzKivC847LmcQ
/VO0mTOdmQ0KDTLPHyOgnj64PT+hva2yxGBhVDIsHIDWsubWHNO7dRefclmDVcqfCwU0sCUlRGtc
+MOMiHuwrSBsRhU+VAJ1DmNPavMyZ1D11wzn4pjwn+g2SJ0EbtyayIhpYcnxAjcltXBEh11U1C5Y
wLObengFWe359F2CTcvHIA8nQGuI2E471EE+K/E9AHJiUz51aI1lm/s+s6Zu3ze9eIzuaAe0tAsu
nbhzY8EssjG7s8xLgiY0w4PdAmDr7sjORpfupmZw/nhwlS7zYHMZo2qCN+ciMa/wIk38Ou5qiIcH
a+0mnb5+K/yPg+P5NW+bFyfeIOksFzrUpl4TUygqVnUb4L8qAfRAWqycvXoKlZOe+OgcwX1YsITP
mjAckLzGubJYQc2OfeCjI6TUhSGU+APKHKYiEM+x13Z7bBoiSxf0BanakE4NruRkqomisgTRf5GJ
qZuYCKV4KbDtPAGuCE75Es5vCjcY/lK2/+3zbNdqJdYohsue4ZOTrHbb/0ywzGiGmljjTKAaApTR
BtppGfhE1f0VZXQo8kXuSQH3ZXcSHp7TgHCsbC7DnY4vNSU0bNqzRlFPy0kSUt78kX6VyJVSdQXs
G3yerNwHHFu1bYSBb8SILi9wmAr5KHqNum8TGFJf2TPQaMSZRzYSKfuZ0kXhdwkaSJz+zw1Z5P7u
58A242lblCKVs8NeIFS0HtUAJ62P+A66UxaT7IkNyDpDebM6190h8M3bG07sSlTEa9NkDya/+Z+y
Bz2TaSROe4S1XeEmN18mNojNxEadztE77ARMVQQI3vaT0+nxsYooAQQ58OfiRfU8jerx14TDVpVg
cLPjuokFmZTtxDdGJ5a4W5k7OOCEW3jf3eXcrpowzxCGjNJBHL92oNtW7guMLXzsMrppqd2laFFl
4uJmcfhPh63QjBvc2jW+UgYlviRRmC5qWYLNtewu3G3lcxhq9bKZEli4oeeV/se9KApD5ch8TGVu
OYMPaPquPx2aO+AdHQAu55v7a6hzPlG+MdGgevkNG0lKOGEC3qkJj4bfPQ/CtwBNmMO8rF53XCqE
oY29PAhdT9L8hQh/lD1OB1neLRJS2xNCD7hDOG3Ps0s0lX5/BZRY2NVxkmaphs+AY3wlSJ6jOnvy
X7r2IippR0erKC7OYsEYvKtMFANkCteSRojXd5uaw3n7GGz5/Wbzs31Tchqc6tk5k/+GxqVQwJjY
h1aZ8CMBjhecXiUlGNOFLgvMNSUriwdaa8zBjknZNfiN0WRyMsu+quG56356UHo5t6EpoAopCTK1
os9KB9xA154d1MK3G1BJfNaeJ8sSNw1+y93QdlSu3ATbkt3CyhIytah4+eDzSzxLCCYIKrJGRRiF
ccuPvcDEYp084eokBRW570aC3i0uqPp/g8wf1dTmy0/922YCk6kq0KQkWXMQFPhvi7ww6TGIZyBi
pIWTIuqunlJCFKJPPuGomkdPi4JRlVc84po2veqGECb2S2WxJGD88X/avrBvxzKV3uYV5voQuSlL
P6qYJEUvDBsmMgoYvSyfsQeWuk2ge3KSsLDxuxtKqCPUa3Le+jDshFm21M31L6fNLR+7oJXKTNLr
KaI79WoRqXCltBUjDVo22KcH8op0GeI3y95Uill9c64OKUo3U0DuzwrAVraqQNFwPyVrE3GmdMSb
YxEI+O7wsIGZfkqJPzUphHAKHLvw+IrKVSqCIXkz54/CkUwAQUuctkdpyPszOMEl+ME3sM1Ptdu3
NO7flJbwnROIiU4JXXtZZWLvLGIgO9VoLZJe3E5r4NxwW9BpV7Sa8O+yjIgVQAJwFhsa3gyi7gL0
d6b8sK1iQSBratuj5gOvzPOjbiV8vMkmurEhf/it3wJWntlr3+YCXzy1xkSWrzwSujZxkjG4JGWN
/210XjuXTkXTHoFexRs7qctI6g10YSHDblGF9goPaJpHljp++7kMujsO7jT2IE0nLswh/w4HcG5F
H+xR2phwRCmveJDJ8NowXfuPwqW6SnmN+WFhZp041qOpXfTqB2j9CdnTb1gKO2lP2/hZ/9Zzhgu8
uIDnsLLiwlpHurFx6Ke16W+k38hqEysW4Mh02z1hhhOL2ww6CEGy0Eb/il/tLglc9uMHHqb67Gob
/Deq7RNDUkXj3UyYgEzMh9PPAg6OQgpdtFWryj4oIdbLn53XH7D/Hj7P7RLZzZPCz3gxip8YI/As
tFjtrbnawV2IDYTfqOMB877XkU4TOCdfflXqAxjZT4CJVCQ3nHxsVudmxWX5NPcO8BcoFBLYODxR
PpGe7ohnHZS+MXmLSxTK7KQjM52FTUUFB6hZgk+S7c7inblF4zw/D47O8QW2XWhI5vWzq9UxnRDC
DLRMzXH1RNMv3xvtZJhHo1BcRI2x2ICstlOZmXWGQAO6TRLO+RXRalRRveYJCD8ESlcYl2vVMAeN
GAmBAtJhMb5sE36wiLGkt1RacSLOxykxlvkJlxZGoVOsS7Lu0aWDodL8OBePcYk1tu1RNsXDxt/0
DfbmQbX6XZe/YsVNpt+yW7KHZrvsEaHUCTk5mfbMG872UaK0883DwUudxQMJ7AkxGpB002npibKu
bTflV/bU+aIWbAZtWREE9J8xX3H1mGAc3iJHkaUtVfYWcJrDOUdklM4XGrPpuruAlnyxxKp9Oe5G
7orJ07EcVbomD8Rwo0kl6Ljo1jKQILw22AFGdCidmuK2WdhaiJ28oBe1SeoqPrUHD3GMP4/DP7UU
XXFAOwV5/h8AwQneOuqBhIE1oa2dMlXdr/WGaWNdAqeWeowJHgQcYw+0HPCjnIKfnllGINOJSCAn
rTJC2nLDYq6+tsSQsPBP6/rtHpv8BVq7FhP3ZkezMKZ2C26bdsvqreHmra+sB86hOQ+tl2h+cmUW
fCfiHrC/keSHzyxHw9O/Z3kK9fP+BOeAFhomHpIFMLkc4jSzxJOgnaa0fOr9I3IFyu3tEoq8S0IH
EJswQKHGEBtiGftyY94OQr6JlblUG1uK2XpGk1i8LKDyCKGNTKefhZYQE2ydw6HPnMASt1S1uxnq
3ZPP2iu5VviPfdnWJWfNUZRpS+jcAPVRJjqBlg9LKe4MrZmov5SEmCdhPaTOpUGlML5rIwRst3ug
JcRpC4zRhr5O14ushQ/WNrof7ie98+o8meFDJV25YfQbTogZPmHzzEGw2qbpeOxxl/XYqS17NCSE
GiSAC38Rg6dqV4UYizl/L7+5MwYaHBfBdBBZOdab+HYSMvksan+7eNycxsJF27IvBoX0qXi4SsU2
J3DfRzSurz/8kpZwxUBbAmwdNmr9f2bTEvVlmhdJ4AKpHYOjJN52E8t0k3dLwsig0BtQICzCdZ1y
5fPenvVDMK0F0XX1TdNxlRxVXcSYe/ITKVthK18X9vKIGw3h2n0o0E2benYN7Wr9vWlI8/yJ2g4V
Ukv0zHmzv7folxCu8zMqQlZ38ZUGsdihp7H2wfFUgtig1VBc3H9iXrxNNl5cUDtBIc+P2RQNgW00
iQetaH1VDQ5m8+IivJspNkYCKojPUALx8hhGUrxAz3b8ThLZIx8j/U7oc8CI9D1pRCMRmRMu9pky
+CjjpqWuAc7+vCAAyjsmqETFxtYcER2DKvuKKWaPzi8wJsez+NqvFVZuUYfaQFEdVfXF7XELjSSO
qN2M5WaMs46xQLPu263QZNEh1SDL5kq5jIk6IY0gpLeJ9/brN/xOoXOPCa4H0aAtKBEF5/1ygiTC
tpg5aIidJnxGIYU5VSfmna/5x98yBIP8sk4Y5QmuPps4YU8deCJIZemhEA65rHCvF9x2cc3WeSZn
/CAWVVxclnjnYC0+3koHyz92l3XbNgjhUo/LN/QnZkvzVW09Hq7ACzx+dcSOCy0o7igS9jltaM+X
LXlPrkJwqKaE+nDvjChMjhl5gIAQHVEUNLwEyiALhmcR3t3ZxlH6HzxX4CR3vxfCkWbcCHLj4drz
Gi/3uiDQ1jaiN5g0RVMvN3WEpgKkfMnYu+Ad1zxi77yuuttuhTHWV42m6kHPEE2O9/JzOY8CR6Sx
slvd4/CCH5t76siaGdTn6YsVxm7Vx1DgdEgGJU5UVS8KEO7ZiQSD8BdQQZce2/XOG8onZVrIB3xc
tujkhrFkBYHEs6UK6tOfVhVf2MhCl/1ms/XJHuRibIPgbGMJBgkeYLnG45ioK+zrn7BbvgT2zvPp
SZ7kEjhQXVZlfN8YaTELc5YAcs/LoHHZ8hpNEH98Fm11nI0bBQFuVAv9eb9g3JFlEHpO02iDH7vm
IJWBmuTs/RtVzBPGunUpp6V+54jo3jHY2iQBtHLdYapG9ykF2zkFGGjB74rCAPH0FsV7ASfwGoMQ
hfxYMG4vLMpTXhWH6ADo3S4D7ECJzd319q5pr+8sQzAKwlF5aIZlCKJ7hKuKW4Db73oCwmCE3yKz
hH7n5LZGwr9yFFkyGn4kva36B8A4dd9KG3qtivJQkD5eeE9KwF7Bkg4yzoaErKt3G6kCKvNLB2fE
Ytn9PN0ql2x8Dc1dxG8F2SXSvAklk5SH0RM0rTvuK7oCDalGjWxsTfExpkmTTigtkuyaZoxFIM/b
RfunM7z00bzyiUXDdj/7BCp10GkiqTwpXe6ELML7c39I/xfWDW7fXS4BHWzvBYCPWCDPnk4TmLTP
xt/XeFdC1j4KFAc3KQCgrBIH/tmnSBALF2d+01Ys6aV55OPM0FJJ/Tzq5eJDhee2RE94ZsWvW/k2
T4GRzPOK9phNk2eLSsmuoDoJzl7uXaiVMKoSW/N2nWC3Udo7dUJy8wAIbJmGCK+mp1OXonIKvXK9
xddaKO5Vv0j48XWOwXO0+Y5Mk9gy5T4GqPX6QzqeIEUu4jSiw9z3d3lQAF4HNrxOVmimQzmHaKGe
ncSsECgtpKnCrXfmThjy28PlBGUGYajWtMWHYgpV6Rt4ps/YxB5SPHiwBrw8K7nkdNiTBGQjt2+3
IA2/WOwkUp4xfXt6tshWjmCrIpPkUL4zKgOwdBb+GtgDUYXgZWf3qn0JNmQ+mkQiTCXLFv8vGBhw
uPzsaNsMHNj4Df9IuGlkOlbhBaliFHmwlknOG3UTNuhXIUhCh+IMTEL/xJHNgnY7l18+FGMmXKEJ
RuDmjgjfyrBetqEDOTKO0x+/qPmdFA5GCIFC8V9oQq9Kd+a047NZTgi9EId/mP5ZVUydQcidL8Hm
qX+1wwAAqwEYTzUK7cLHdHvWz0pcc7krbbWltjYt00dmRzJOK8jd/pDqVwch/M1U0LNBMcmvCmGT
babfb0Ynj9OyAcrxgbbyefRlrjcsJ+0VmEvqXDSuismsFn4WJqPdMKW8uM8DYx5zLS15xPgEjcWt
kBkw/AtIc/lLXLZRuuqkhN51fOhxHsJxoYfoc93riLumZDeyrZtdemXwuFUPetSxZEKZ8USV9aVX
JDzGxOHHZK1T3QzLh8CygpwmkmhBUe5XjVulDl3EiglrOOYmjLg3SXDawqpUAFqEfChho5jogLjV
VTeVjPbvVRGWRlsLtCxw6P0oo1+acR4ykTvF3RL5pKicGb8Yx+eWiicMW5jEAwRZDGwOrLWrsswo
pV/laBdIBKc5ndRmejgHMZb3e/Bzng98Ss11BuYdT+ns7iVZAuEefZMKG6vGdK+g1BAmnfmNkD/Z
y/Ao48Iok/kMGzE3tZIKADjGnt3BfuGvWMb3neSkaZH1NSjtFxl8WcTwaYku06ytqkBxYYc4UYh+
hWjm8D8hvQvAMFV2WnaXTtBd02Bxhb1SIBvo/tOEUHXMJkIEJKFM98ZKl1ypbWv7aQJhggVsgWLv
w6LpEi4W43Pgu0Rb0Kdi4PYY/muo5ZuTmrNxK29w+FrmsWufZx1MaMuwZQ+kEP1Undle2+/dQzwd
en37MASqASTaAjTCdd4eTNSDmByY0/NojCqxdomYxzQevFQUMGrihisBNd/sWw3YIm32AETwMffO
3j+L+ajxr9VgyA3gbNg+I/uu0uiCLebmHgsKhSSZokoNEpIy27/nFCnE39UB6ezlj1JaKMTz9to0
vYGXXSU9p8DHdHQlS17OaDWadCDW5RIxlXtBihyusni+4xGrveZujkHfrlIsjzpLtZp4YdNouJgm
sOmyil1nNyA/sncCEnA23pq0/zmK2KLIBmkuB7QxGmPEyeFXMXMJYyQZwRLibglNbhZCZW/ZwwGT
LKNuWQpW+0GOP8xOoPkwy51dkTOh1dDndQ2DceFKLOdXbZjQEyjqmNHoECxjAY1DI52Ziwl1x/Nx
7tUNfqMmJO56zrcLK9WQXAQOUvOg/+pzfgRPv5OFjGeHV4oENvo8cZqktp0Fr0K2qh0NbDGb2vds
r6BJjedZPURn/NNhyDOjV/psUbeLnbPZ9q+JwgGN2C+uHNd8SQSYyGKsqm2q/P3zp0QGhNeZ0YBt
7vss1GJRTSn7FiGCUyDf0IAkXcaFffPOnzQXzliOvF+jFNN7w+N3TodPqGSyT+IJ/iTVrNo674N+
MIcN2DR6xlCuFDkYx8UxgMtHdmcQ1M0RMUQ66MxVxb+ul5ymN3f6szOMHVQYCznKpwsrMf4dfKAu
v/WrMzb7dg2/0ki156lrqxScLljDUJQrbblhLc+t+f1YJS3y25PbuTvECqg4wOaUJdUEP/jA/76h
KbfGQDsPnVw+gAYWPtYf04j//iVnDH76adxsF8johlmCEiOQMGUtRJiFQ/BsEukuv0fhkH+PQlca
6a45bzoKhkPkHzpoXSRh2YbSRWMEOuE21JGNUTtyEGgqF/yuDVw7dZszU6P4u31MT9VAHnlaYRs1
HPGLnCTZQIjMaIAuacDOhXJEKEMcVUy97Xiv7jOr8Evw56oVY/XYu4sc1dNUyc+PzmAyb6CFquTt
cM2ZHufG52xcLYza1nbxh0Rman2ciCIxwmj4MJkML7id52obS6BRoiCPgKluSCBqmnYpw7JICfTU
ruKtjK879C4BH+z+Djz5gCqpliTnzQvFOM6P2NDvqgWsz59l1YQlrA88Hnj7ScV+8In9Y9ZuLk49
xr08K6d6QhUpGfXBg0ONfHtvO3JGoCGc3SgGZnXtOGw/TBqSjCuGOJxV85UFWUY3hO+WmTQK83wd
6unLjyfjw0uRVEL0HXHxA2VEptlc+LvncPDOTDtLdrh8L2w9xPOcHYptoZOa4xDumMhI0WWzR62W
E4eib9Bj2Cn5/pPKo8EniMiPZdu8PU6lozqU3WdBtByIE7fIwNtg1LV3rhoGf5MpICwtDbQ9V61h
StRgHEjZn9SWh1ZOBUAIqQpKFIBxvIr5intiTsRXPs1Sesf2Gt9MG/pGxdyP+b51u6UZRVieKgit
XNcissf8Ic9W/TeZnOUX7SG2l/dYhB4pyUpbUESqHo32P+6H4qGH9rQUApDwqlTVnF9e5XCO/Ukh
aTdASOH8DN8ci/UJ6VTPRNryJuozsJ8PcMbJW8qVqwkMjl2bqNA1io+SdTW6S6bjTI5AMf90bTIa
R0yUGhg0qew5wGOgxzKrs37slWAm96s/4fKjJ6S6drFKCSxp75WyvYtdqgX5/xhzosQnyNwVM+df
laeIo+0BFQ1N9DFwSbzLtKR79wS+ig+rmrtgRjla3U6Ctw/V2ZeDHbvAsofP6qpWLagfYOUJzm4B
IHhyJMYEXI8LJM4bpuWKfo7S9rQ9FfhzBg0RDf9XhgmxVFQ2Bt+UnkKwYzNiNdOtAB+ZFklo9m8F
pTIQXKks1jzCwVGHfkd7fkyZA42w3d4ZWF7Pp3ENZKND3eQ8P9wHrQE7IIR9Z1VeEibnVC2Z5CHz
KwdwhIxh+jhgqAv0PlznTjWmw3PzpZhdQm8dISR6t73OvYo0hLov04sX7Hu1lt9W1kpAkM4vTwOJ
9luEwhKlfIbxtqR0o+Cuwa3VLWtUNn67Bz2iujgg17S2qqSZnbk/tbisFyJQ94uzAjrCWJY8W93C
qDBU/1W+U8DFiPvHsbMJS8Bzj2ejoLVZTNTVs3AtfPDjQjJZV9Bi4tE2zLWZ31Uxjk597rBkXL1B
SMmvl1N/JaUdOuNByNHqANbIrLw8OkQCw+u89nJ/LiAIkSkwDhVpaEUli98LBhGLD+Kd+xThwU6H
E2jhYT+/tP3unEws45MAx2fPELEUus7yTc6d/U0znWLsVx2SFa5NkQk+TDG+g3V9XqzyMTLZDREP
Sq4zprhR3O+YI6gAGnOsWsruSq4unDLRqugsyva7nIxCR1gVtYAUa7/B0AQtDd8i08XPVJFeZBsb
lAFlWfHFRj3VLNNHOHkgJfvWuwLR4m6+v6M7xpPD9nBxtmgDUgOIsbVyo3d7rtx3xIRnP7DNFPr9
9UhkxloGK63wmaiDEtJg55ftILY9E1DnXv/pk2B99BBwB0Wm868L4nTjbhh3PHIt0Mui+76BEIGd
SnvrdOiEocqPtFHjzWukYX4XEp78gyu5mxIXfaM91qrVumXVMTU+g9Nojmw5uPLAGXM8Tj227JpN
4bjJrjvld3jZq1cy9rJDqoUuk59IMEoMfFcmaTPSdK1JvbWcvJM8f2ye9NL8xgU/cL1rxrrRoqPl
9ysvNUoxxZWdRujO6HJMgv1ds/JwOB8dSwXWz0G9SRzdpQyyqgo99keY3WR9KvTL9mImdY22StiJ
t67GORAEGyqRzEPkCTWEIex8pYTSpYbVSZzbKpaXxV2Y6GY6naPJHcYvCAmoudynUU8k0FfufMiw
GGi+Q1qXMcJYHIs/HBwPG7aPFozsnFHzHLA0WoUn+uxDu858sZQMQALbzmc+DR9IBmo9sGspdsiK
SBzfLOAav6dB5qT7tSVwAqWMfx38UKvQM+AgNjAdTofGYmKcK5JL1KbnyjMoOv+rVTFyYrQKTq4w
Q+a4HgwYB1lXLdLPZZlDjwPNdFuCbgQ5QNYPJ5HT2c6+CtSkG8zuOBEjYa8RTBS7MU8N+PUsx3DE
Hgk8RTMoq1NxjTkfyoLxPb9EfoHYzXqBgDtCvzeeNh6v7HMqPr9ybh8aVv2sGg5eQLHrmftGYGTf
TVB39SJXYruruABp7eJM19RrX7PXRue4acbt1OJdG3YBfwkNsudqdfwI6SaT+X69jz/FmpEwB53p
I6HgGQry1UMKMlzpOD3A1VP7Wvjs2SURUgNZ35797szu4RRK9QrPfTYlrS2bprikCPHn99GmFZfB
yEsM2kMcr+XsF4DeffIoqZuh2oKL9yS0Gkf0ojtoh1igaN1cprlfoHKMAZHqz80ux8TZ3GWrGXiX
kX0v6woDQFOAxsXtKQrLZXHsCoRZXAdrpK3yvsbBGmD6KJiwc+Drcdqv7nY4L/6otdv/A8XX+CVx
H+Gm1dSi/95HLdDLCZM3fZwTRNEbivJCCwV8M3NOQNDR0Owz2QzgbA/2geXlk2MVsJRqxSrwGi+P
XLBDiokmGfixfZeqEP6LwfxaWic5eLLYFCkxy6nnnq7N52nShI1GoeDaB7QWQijZARfZEV8cbClZ
9wa6T4xkGySqeeuveqOos6EP3+AhqmYcE1NnIleK/nz6OWpgmqTmMnXbjCxq57Xkk9wBXR9ke3be
4aMiUaXuCBUKI+JmkP/jbQd6yyAG/8VPTZbF3EUte/ZCaOXJqpqAi1Lkjk9sN7QBP9iX8PguJ0ac
ejjL7O6HOxAh30JI/qlbNupjjVVa04aTRrqleEfQ7p3JaVLQH2eyAF67WCOItDgktIE4yAh3j6qR
cLm9TRXsroY9Ddse0Q7/djgjf4//gWY6p+A8ur/UYb9yAsz6Dj0cUqauX4vs6NLiJRq/l1jGr8Bo
qUuvQ6oRSHehBElfdMcKQwqosk4UVoNQXqIepvtI7ROsPWK7CAePWgdKU5PzCCfTKSsGcNQaJarZ
Zwjp85MWZvmMcBDnleeK35DwEEvhm3PvjJ+L6kM3FXJQ18ikrBTughKJN9QLKyBLcfJJ5K4Qe0Mq
JKRcjRbULbvpdSHeJ1HrKaPLQzqISW8mGYlTSi/+2UlZAsPwxpSZAaUNKsPQ876MTdHwcHVPvwiM
NEEg6ow0vLcEAry0jvnQiEBLYVtOhtfJtQz6H08ika/Uix1/dR3R2jmwrhgxAiWZ4woOG5RF0Ug+
2tux9iw+FtoC/NrmvYmIBEepnZdBLgKGb7pfamPuYlnnreKLQ36r3mw6P4s5Z99fhPK8Kr6vFnP4
1prG7DIm4j8nYlsqdal6ZpJzZIzPDdv51d5Q2Q1hqOv9Gtj0Rd9jGpUol1dSo56nveapMOMDY3qS
tku6dAl0rzSkBevIL7Y/935gs14AIMlIbfZDDgkI3rjO0zx03sduyk/m0US2eZUeC664aQwRqbuY
gT+4sFwYlUsX1qFum8DdooXUfW9FCBIhmoVP99EhvV+syGSJVEuhFAXOo7H2HTDvYNeOxZ4PRcS3
ec/sVrDyLAt6ZeMMJ3dKkvXP+WO0lqYumJrbHZDYbx7r+OzHIXT11ihvtT4jv6QuzuplRsl14fk6
yMjMSkdH6c8t2RUCqIRszAhse4udZvqLUzS+nhXLmqr+T0R0gbbYcpf8ZQJU8ThKbVd+6Cw5sSY7
nKZ2VGMwuXiGoKWpyCw98QZoy4htP2iG61vPtzODYdSGXcR1a2nMgutwlXT8saDpo1aUvwGFqIb1
dOp3wSH9bySVF2GqDTwQ7gKDnQspEGfsi4SZslcJR7On/BxieuFAE3/IW8YOU7SgiH9IQr+r0ZhR
yW0BVuCYrUJz+PHL4p/vrTRniQDCpZpPNzFcmlhhIFF2KjX7hjzUixjkpdB7HcjVOTiZX4Fjs5Jw
glNbXaedOhwjhYXQipqmP1jgwyoJ8hqPFKvcSZ7HoE6I5E9pJ/fmPjZJJGTp3dzc+pryW9GgaLZO
WtnBYBhvVjVAxALxQF6ZihsX+Jnvaf/2+ByNkNMLMdn1piEqqN0rLbtkhRDntzQEXByKwMnyxrWZ
iFJGYbxsCricyeabwqj319raIpy+hWfe/+pkwgIz3pC6hhc4VoHcDlKz1oG6GgmWibCYaqvxEkKN
6MccRWziyae8VWKI3OypZhyR5tgXM3nkeb/+aenrVW49x9JPvC3p0CvQjaovxJ+cCZMwE3b7mhC6
zxcZR7SPtFGIgyww96gapJITNtiUU4yCV6xQK9kc0uotcXFj6FhcrcsXxsAgv9RzzY2X9GmxJ8YI
SvwfHOv0FPcvYGxPg3Ccfd87J7mpk0l5BzKkB09U0CPyyyBz4zZh463AFRhvrcMnV7xn7LZxhUBn
9NWmUmyWws+3v6U+aLw7K3+7ZLfLqMMLAnaA/Q82Ep6oI7hftUuCKZEnDEZxl2baugkmlOB8ipTa
233y7WG0GDJPDz6YCPpTmmbNbw2V7rIcdMgEnqdwkcteIhd0W2YzuBWt6xDyeWtV1tezHF/sIAmA
8eImY//kUUBcaFGoxufb7cLrxK/w8+T8n3+xq7UbqYKQ4EfNsMoOrh4wQOhLiv+MJBRs6bUDuliK
0oYcayCoblq1J5TWEiRQYu3esUF5ePp3PZvcRD3rZYAXxZZoQOSYpyfG3BI9igdZv7nnT6RKbx0E
5cdoXY49EmDSes0il+7UNDknE4lzVbg6khlizrwCxUptN4NNBbOnlNA+2g4qmgZlSO+zXyTSlZW2
F1wgGUxg18/OOqZzJxeuikaacLeR1V1gghTze5wzzaaO0X+oeIMFaK9JP0yLDQzP3JjsVRtOyHA5
J3tOh7WFbjB804Hie7ehProayJ2SH6ggUana2Oy3BPasZj4EsjkccCe6qVSiLvMrOmLNKexW4huH
pbDB0Cg7BKOAv4pCh7H0e5BElv0xSBhYmN1OMm091yGevAD78G0ZycnxYnV80yYq6Q5lBymyKFtD
zt288C9uk7w0JOczwO+N0HshqWTYWwCier6rY/vqsVMBLknKFZprp561snQ876qVQJQMkoHTZZrC
2T0YjmBCEKgDQdcYxbdElhi8bbSJD/1fyxrWO9hlMkRsf9QifuvjXZ1xby8Q2Pm0rxFMMn0dNgpA
8Oe+Y0hmvEpR41r2KRpBdOTRkoZrD5L5QmmDjNqLugLlJoKr2Jw/fs18AV8406oU6Xp7BmtZZfbD
6IrGPCh39tzWlkAcpK2NRfXYSlyZUKQJsBNpAT+lxZMGikE2uw2WDdfXmon1/ebTuWBPxTkPkiSZ
XroMXAp+4s++q/0PBaUw7+vzZEmwVEFOca9uDHk6ubtwSK/uJk4p9e7wqknzwjufl4xQjUtvVZWC
g6eb91lOXNB9JRztqc6c7CYfMZyw6fVwqrOyNxjMOSONrwBjyWZAeheW//fWDBQq85xUGdGDdtyw
6wCmpHydKIyjsj4wPTLCW5XqUuyDhbBuENTO1EUksRcXduQvwhYZY5T6+T8LWNvYGNMwEZpv+JQO
uV9kaJZBptGhAoNPhT74Tds7JiTdyDQCsD/bqCT672DrUbwhvyrrehJTiBbDrpPUesSvbxfJSYXd
f9E/eaBlMTTVr6slpQf2DNT22izmU8nXbfS+7BT8XkoGofQ4Y0t4OkNbOaIXKEbPB5/GwEnkyLNb
CK1Z4FgZntP+cEnn5yDeruFzktOM3hKKZ9DoZOMsrJsV3IzXiWQiMYI+NnErAZzygnL5gsd10hAd
NhvrF18iWNcLUt0F3ACoY/CQRuPSNjtS6Hrfz0YWKfwJJO/tvx6bcuCOrSMk6m9uzAmxr3HHuzZg
+fwfVPq3q+A/Q7OLyefWeXA+ewW7ofVSgcwt1gdmpW3EQVzmzD0YP4ebgSn+m1iyuaQkm8d26QU9
ueJQNbUhyi8fdtG2/BNO73D2J5BlOSLmidPeqGJLZkKdEOab46H+RCLnTnzpaUoZc/en4VBDpoe3
onYBnycKrNdmg8NV+QivAa3010otrS3MYyY5+8LQGNyJQTtoxoYk2cPU77QlddvnMSxqMRu2789k
t3TURpOlEQRySAtrcVstCz9rikG8I6K71e5eUg108TPyBC/d8U3yJnZ47RVIReCNHX9QAeVuE3dw
+px48P3INknWCcakSlHYKBO1x2R3qO3lpwoZxkQsgVaSwv76GmEXUEcJDDgiE68ieKUMtRlRzo2Q
ZnEf4utywTZ7Kt5yy4x7PAKX98PY7Pek+CXZOM0ZrW+c8Gw7i8G4zsICbFF17aloe0JIXKz1zZSd
laJ3Y49TpacCrjdotGZWj/9fmvVY74cO925y9kZZ72ZIkllBV0Iv6w4WzTEMNcH/2URNP9FlGoI1
QWU3u/HtGE6pb7pdFRh09nPQbCrZpW7piLXWyFUWhz27IEqL87QZSqzqAdXEx07c+bURsb6F2/ON
dZhyFF9iKfwQNKa/w/N2GNnmOWoTji6dUO1LL2P9jFHUkfW1eLgcuELRzOTWRYmRIUk4jXF+qwLa
FspGkQ51ojSV3OgTiNyUrzK2n4lXIvrOKktf/BeKbJfrpp8VcborowlrAFqFMvCvdGI4exUbYeEl
8LyKVIIeicr8kTFiRcwpJZxfmGqoZ1dqdZGSq6U0gYB/xD8qSvUVHZ2hpotm8uHM10pG/1QzlcaB
sqnINrg0bxsz6EJhVAoVqyteo2PyW15Sqq2BSYXFB/oBar6O5+hWsZkh/dxpeblfb/kz7Os3fsNa
RErtpCSCfh61IWRyGNGLVkqY2Qmiy5s27np6+6LPyTOC8px4IUMdd1msGuYlVdoGgFJBAdLIzYL1
oJtXDtzk7+WWJmbDmwrk9GI5l9lmJs5/WNjsaxAJ3eVz/cWuWrBAypbW+SCOchoOOWrV31LUMbwR
EiByL6cC2DgMJi9lvaO76JziOjld6bsUSPNygvU5RqeiYDUfU4goWFn3GmQdErWn5GIwkXyBfniy
YRKtSbP2VTXODUuwFN3smoBlLa+BOndbH5hLT9VbztWis9qQcDjyCDPYp5tKdHlwX247iMwJ++uO
4t1/dafwLXK+IzuEAl598bTDdkKAWlel7aX5OPNtfchst6NqZdvmW7zzo0qumdzIvlJUmgqDHrw6
xBgnIQZvmqZOMvoYMlInSDVZJEf2vJfPb5Nit85q0LJ9aOIVvUGxbJBird8MWPOezNjMQtohFByJ
q+tHrw0ogehQEeDbB87eJxxFHJgW/t/WYePmRdafUwZHOFemeFIoAz5JuxzyA0qqhbmKEOg7PC+A
SQq7JwN35UyYXtlvOgz6q/mtsEvf0ejLn+6sfIfw/y1gDMez76wAPqLzTGyacOA1M1pYjhqXTfV2
pM47D4YMmq7MPDat0qqvwFRG2Mw45ZuzQ98wL4PlnkV6bAxu3DQs0HF0MyqYRLC8owAWavTN9sia
YFqH9zagvB9zk9LgL/qir0volyx2RuTns9A84CTtYeLC2F4CuBWJuWk945kedMefBo2l2Bopm4Ag
SU19UWvlKJRuZ4oR2rNZrvWj8N81COg12ZUzJoFKlT7heezEEB7iIQ/JPPBS9SYM529bH7AAXryZ
oXJi7upYJRUCrvGZ98iYJPYCKCqh8IaS1T0Es3d4UohKWYvLXRJ5w6L3WY9o4cpNpR20UtFH6Iym
u4KBcAu8FV8O6g9zytwBfZrlzPDNHrwpSstZMbL6T8uSHczWYBdKv0f4BqUY0dN5x+0NHdwkEwwx
K/MEFiLEZM8o7wjEb1eKsoHkvGzZKZMHrwr6GTxww+57+nJftqCmfi4ktlS9DuSd4I8PAy6ghrmc
Xjzt1RKX6/QOuzUg4R8X8Nv6WHnsTT6Yd2Ayi5oxxvlivotZEqo+smkirh8z9dXCxplj+vY4o9ez
LvAzQqt1Qh8FPPvAXOqB7OEGkgsQi2UF/7pf2ZW5Uyx0FmETkEeoCkGQlh8rY0UmRuF/0600wRNC
tI0TQFE2TUgmTaORquz9tcB4LongcDxMXzOKrfYuCwLhEEw1y3CWTpGahHdYk1EaTvNRfnqGdnrX
WseSTSyZC4D9Uk3wcT8W9WH1w90GYvuYlXTZQ+MVcfr+FzswL7EE4g4jJhTgxwTp9Bb1Exss+Lbe
+T/vtWosfmjl94yemj9GWGrGyLfeuzoL2UxT0Ze/KwrNQVLLFOcUsyQYhMW0STHFcCd19OCKtzt0
OAaDesjtMFOvFr4VkTKg+PbiGBLGM9Ip1Etvtodl+zaRUfTsSTkXIOvC+rXFrT4uShrZ9qO2VsHf
q7SiSt9jyZV2Ey6mTIlLWoULlNUOTrbOoTXyFbSgo4ect6QOogm2HaAoXisCUW9Nasvh7KhTXDko
2545SuuAq31YUzBZDEiiChHLGVW3ZUKBsCcqYVLx17cZy0lIjVLTkWj2PEHI4LT3SKv6OEe8ke30
6jYti6oyDNfWEJUYviR751s+OoZedHvPoH3R3Dxf/fdCgTVy0yCGsElqNa1C6V8tFkdNWo4/rC5J
g95Qr2sEYrtFN0+13tqu0+NAvkXAt6kVpD/e2diEXWZAZbky3SggZxHOYa3jbEgVNSv9E0ICc7hc
NYj3a/zfnpiN7AqO6WkEm0XHOc4s244zGLx2u2Z6PI6iJfCQJWw7V7BUW8xrqEpkDG1tw6Z5l5+P
cDHb2UvfVcKzOZ9mDP60v56KRpIUZJxmH0w5lth5CI+qh3OaeNLuyZNx0d9vmRUbHW41h/9zTduP
RRgiZz4K/Y7sNK0jTVoeIVorgxxfI0C9w3Y9go6RZt7u5BjNM4PhUUURTsN6Szm94JH51JhfeY4p
TPLVH7McktT1ITuNMST6BzqUP8HTj6CVYe7QP2+ps1EohZANJkR1IbXICSxX9fOAJHM6KvPhhyoO
sEIXruF7DNNRZvNUdjLy+T7P9UCuX2G6jVaygacezZcDLF55kpciRgifW69BBhNCTMkP41TIzcd9
QmvzfqMvAy4NysaztzD+XSUYFQyjUWp6G0p0xwcwF3yGNnnvyj58tHBhwxeGpRTbp7LtfEQxenND
9wDjOigJoJ0QxqZxaHPSkqNkJeIZ3ObudXrFkb08aSJ//UpySkWzQI46HmEG50c9Fno/Q4O7uBCm
sAeoZx/lwI9aBRjv+87SURPQzOE/3zhs2RI13gDdR6aacIavDWJUgV8WkLQ81akDw9Zg0s0KeyzN
OOdvcF/CqAgcTkVbu3dXPxROdLsyaN/oaJsJ3OpNVwtd4Wn0G9sZMvTbhzKGCsSyVfMrbOQRC0+A
lJai73+kmdZ0hG9o7t/jbzZyCJ+/N3TwZYvir475Bk4WtnGn4tpQXmR0bXshk+rtmPgAs0MPA+oE
MQlcTXMF9hNU9zS1tV/TOvFOOiqh1IqOyfYYWUNHEPX5jKjUenHESXNoPc/mVQSfVKaloFSD8F6e
f0hOLQjoiJ0/0lwWbx+oJSOkE1O7YX98KfErtBGjj3leoho0MM5jGaqZpgxW+EVKNZP8/1M8P7B4
Ro98oDqEPpkU3rXy9LtiQpctKCJCDoGQkYqlOZBaq4WNx/0MYrRtJERbLZABEonFqFjs84rOFUe2
ZMnosDR+dWkbkc+ZXZFkaSbrWMl0fZ/fVVorRRCt6deDlZyj6a7O3L9tEn9W7rA5QOqvrmGPhxht
b/fYgIt+6VpdwsbdpEq/SdxiBz2XcHqppG1EwkbB075rBUZXA4JF+eX/k0kDqzM4TXMKtK+gefGM
sKVTJQx4ls8c8b0tK3QQ8dk1SXGRcDCJ1kemLt9Kg9SiWxbFSWb9WZYm40SGL1tNYMiCEuyNFlXQ
sXc4xSp95SzGJMilC5TYYyknH2dOE2vfnA957njh2KQ2kQGTj4UYm0MZKzigVENp9xSuH8eqZ5Ie
zmw1aSxGRAxBpN3Z5DNM1/8wOH1tI8ZDcD7ljTLvzlXY827N1mvwaHQbfS+vHj8wkNtLJr2An31s
34LFw47rwsrugpp3VKz0Dfya0HckJOgX8O7idylZidHZKdhBeQthPv9W3mm9TwPkHDqRq8p7O9aA
Qc3K0XFjPTLV4HsNnZ1fwREIYq0wXaVtvQahDqaasKSPqqNeuriq8EFzogV4RFJD0APr4y4DImdJ
Gz4YEnEW0qESn2ESOTEjqR4Fe8diKcYG9GO5qO9XJh4Z/pp49pHmb6irCMIrWVhL00YWlxuAK6Oc
7XsTeCdwPLBBki0IOIPG2ejWvRJeYXh1/aL8/aG+ukv4KuPcwcuAeMVDi6nYD4dhkoLMe5RCj6II
3ltCd6Xa9bFJzjuD8xongDZjH1GoRvKsBboP7NyJ7d/0wCOETEYCFOM237inHymUkgRUSBKGgUsm
8kva3hrIEiePQqSfxacJ8U50d+ejKMdHFDahTKCRJfgKPehp45yJi00QGPInsRFyf49iy/of6RnC
H+au+docDaSOxxBQDAu//7iUCsn5Vcl8RJvGMwwYR3iN8/UQN2kJHTINcEDB5WytCkQlIKgRD1mI
LjRQi+uBSvpWtPVSjkSyDSL4KpyVfxSO87LlXREG5f2tuFR6+MK7ppjRty4QtKVt/3tB8BUSbkaZ
tX4Y6b5IzT2wACXmF0CCzhEuCGCaB1Md2Ga17HyCYFxA3M08E+pakymXIT/lEKwcJrG5I0kwvOLU
OO9hs1zi13+ImjbyTWRI4KZRuKAX+oST10WZ6H5HcfkwvTbDTmYjI/63AqvD4Q306wCKMprATYM0
SNOLJzdHxXbLRK+iShbX+3ofP77Iqz1AI9W+zQgYn44t+O+Hn9jK2AiPFn9iIz893V4jmFCu6hP4
0QIQPzniaT7qtgxonoujFagjiy8PaloD4RH7p2MFBBSBmaaLVrkAtuwPACRpNQ7g6EmfnFBEjhLJ
rUmmd77SgNJ55Gs6bcuz3ouPgFFvfu5Do4WJ7/YSLNbHSmERNTgHV46ONqlNEFtlHNk4sYKVusxJ
xkdHn7q19Xxg96iNirz2s85xDyAmqquqamtiQSClx5dDFWXl7LykO76lJ2FtPf7mbsNckzxsxrQo
1UnbRcjOl0le10XMgt+dMneQ/Oqoo/0QFMrINzPPY4wfmM758AYKrLAkWmDdk7AIAFJFM5z/kFQm
Guo5mHVW+fbSLMVKGCdFlhANCcmFf9sPu4iCccYGy2gEauoujtp1EpSWDsCzomHT8vVQZnYYDQ9j
Gj8bsIUivNaI4QW3MXnw6GYewlxHnZsX1NoyOga/5RLqFUram3wrJyWJS40lXjraYIQZ4jL9iide
6Pkt+n/228C1jfjMtlsywmjmsnKlITwc7HwB80WAHMkv7gtRjLHgspx5VeTxVio10Qs4QHcvCf/q
mTiLotg9qslTMCO/EjghD8QshgVOcBxWz9Fc/k2ROoz0bCClGsGyuTTq0Ljzb4RR+h0SDHVv5PTp
Dg+Xq3pPHw+81w7Bd7QxRQk9QNMjzSNQjYYgN4UOXwzGdOguEcc2fgJb6YNlGdCw4nsv3dRFAJBz
HieQidNl30AFCtANIWuOFucQoL6n0RKJOrG4vYtnxsHrkFvBzNoTIg/aLDDCAKqDeVfITzmR0tjV
+CZx8j+u2x5cIDspuJKXJlLmaAdRjcmkn0LjrnFJFpvlo95762NjaAwOKoYI5DFunqZjSB4sg3Xy
+YZb61qoAM7eGXhjrnwE9PIhttlp/L0e3Bqemb3nRcXKG9wABRsiRCivvPPXfVAjm0xfkJvhH3ua
l6YbKxHLyksCarhmR1qxVyNRYafaShnV0fWE4kJBjwZ5uQ1APmV67AB8VkoE0NGuPwmi7Y8B+w7a
bW7FMlA9tfdlvjizEZFbLo3Edk9a0LnGzqQwE7nqR3V/Yb9byUuhhE9JgTCDP3hf4PzEKbXst+V5
Q0IUJ8+o2A4ckg/dEJQm5ahh6uoBH5C1CP483Kq8BqoSuAvPonwHTOmLl8DhJWk76lhJRnqnN0uy
ASuugpbfVZ44HZ3fbuywozAOmMzldNCZR7muDcxFM7rIe0Fu28YQjAETRaacHsdkiLIHl/6qJZDU
r8B20ns/+rRE5SKcA9D7O6nmoaIb/4hoSIyXZX8FWWPFckNaGzs0u5oaf7Xz9RTHlcSM2XNlaKAj
S5UMi4VEM5xiGAehGAP+yE29r0hHJ9hDXKWaScjMH2v444rBHpJGNKf6bW0l9+Bbh2XJTm2iF1ZA
uVJGrQ609NH55mpxJC46VRMZlMwkPyZ7Thr+c6sLJ7uQjFsOtu+peH5476ZnkDYMdvb4STqxS7gV
2GSA3lS36625KPDp2vAD8CfAA47jmvXrXj6BlDzPVvXAahTw3sbr4/+uqH/1PJPwgs4wZuDbHGPe
g3qOFzzJt8xSTnjUYA0Ywxk6Ssqs6wLUw0IAGniMviBhzOa3RsvXGaUhLrjHsjWhaIOknOeJsMje
bqVSDtFoLTM2MF8tU90yibbXilhR9OZh63Po5W/EMUkg1+0G3gRvZsreOPGli8kt5w/QEuWyK7+J
egdN4U6UmGWsK2UltSTAxPoUMY56FT4dqV1Ik/t7QNQJprexaWZjGTcbHKKcl1jGXVBA18FCwoCX
l+8wRkXMrHjnKXbTyg+Rwn2YM671TqlhkVmt8sabtUMaqGQIx+1n5zGv5wkSt0+MaBFAHEFbYa+z
0kATBGSWuV8HJfBtZ7l6+dgJn/4AKtCkpPxbtfyIfP79xjyCdDCI5Bf5Y1uufZlbDoFzlVnLHjar
jCUx967PMaeawNQO1++LJXjtqz1TK/4HfwpPPwFPMfXaxQ78VNagGgHfBOKk5zaa36It6yVWbXfS
Ve2q9OJcu8SCbgC7P3U53DoywgF590qmQNJyDinEro2YrVI6C4mtRge7cm3AdufPPf8P14yTMYSY
u/6fIsGUXPGdGMvQNVgKMvof8JFPun37mycJqctkLMc/qjz2lm627UWVfPrvDs8MjDc0vQlyISyF
je7IOSfNNedMDoHFjQT6ZRmJ5UYIhbdjdvOjpU3SUkkZSrjADO/YcfBWFt8xdOknOrtcvq63Hnso
Y87SLJbECdpAuHbOi5AgrUWZ1hgAx+WX2CR2JQwQfxN7gwm+x0Z655b1M7pL2valReqzAX0j20x9
HdBE3DaCxCDBWROBnNvvEOJac1TxpttCG/AX+zdUupI1Y09H2005HjqkF3s9hS3QIy1IEyhIU7Et
IcaAyn5oFjxeYnHf6pkwHdopIial1l24yD00HKf9jXyHoGXaJMe8HmVmyp/J6BBbNDUMePakCu+A
b03Dg4AoSXegLRC9+e7KE2EZHZJ/wjDyYa+KhauTsYjKVuOwqRhu+jrq/Oy3EkYOcZbrSAyQaHfV
BEQBS1ce4IsnYIJvmAjkR4PCK+Rtxdee3i7PizNRvKCNRV5FKOugtgqOYtpwpX+C7+e4ZY4V0xrI
evaP+WF/Kb/MHF7S/BqEah701S/8zZPDDGh0cWrgOeYmG/hQdUcocJJFiOhNoEeleDn5z1p4l606
GkXP7PUfuYA7e8Knayeb2HgJsNLBfEs7Lt6QewP43Iesh5XfgpKzRSkdbJ3EvjZ4bNpkiTRYKR1w
iTyl4HTmfyMAC2QJ5CiCX6nJzgDzOVRJvVWLp2RwgoXqLl8iG3tMcgvXmtXNpe91apP3S7njVgvP
pPTz4Anrm59kieMUzWyQT3nFSZctlo5e6lnn319Kz16V6YrQD1zM0nxBSlAMp9Q9WofKM7vVMF/m
LJpxJ7ydy9TCxmwsbBo9ASdoxmYA2T83xF+1/qwOJlhdaJZ/CN80vX++LBur10z+pDxEueEUqdOw
OoQyNdBOreSZYpTuaQ3mz57O/V+OK0QZs6A/9GaBNszC39GetI9HNPzbE2iR99+naEWdvdFjWaLe
CDEeMnQ/dVpAS/uvNID96TeRdq2APah9qiq0XJ3HbblZZzWZtnfPFxM2uudP5iSi0oDqsx/Haziq
yPccq3lqk8rglA8YD9mPVqRCQDrfVjhB3mDm+ckuRdjxwlEEExqSwnkJ8wY7TFcN5Wlqa36zu9RG
utMBAUTub0WB4TiD4szutZPqvMDjy7xzZLuOpap9hKuvlG+3Uf1TwyPYxFrO8ER1eyH5fnnelKna
gV7PJR9JiVoPnTjTsI9OI9ST5jaedsBp2z6Iv2g920WWVSvr8YU8xfFApjxMVeG5Gh/IT5zkAonJ
e64ATSpll90xkCMJRxB1RuEtyOz3qF/B2vHZPsRmM8HPvu2qVtzjjFuoDvYXTuAUBHNQJLfi4yWV
SVF9D6tdGQk0TFPIATUnIAtwthrRsD+gDzmc2miFIom5OZPZFnUJu7KU6W9INMKE/aaHXRtWLX97
NBoRTDEiBqWz6dIaed7GVHtuUN8FdQ1q3KPID7ltZ31a49GK+bgqaQ2t/NfO0VxBUb37MvCxa486
oLLJP5wh7/Ts248VgWc9gyaRGECyZuOeO1GaXmfmXtyfue1jWPUTDELcNz2ULCarWNJfZ70qV/kY
sGusmt8SWq27OiBXIcQHLj47zkfUFbfw8/gstJonEQSPBHy6oEzfryNYFFGrAFHKqotjTmB6vk1v
cEPj2IEo5BE7LCsqqumbsc+zXXcne9lesZpbt3shxMZ5UgnAcFAZmgKQrYOOxVAKj/6QMFUGr2fN
tAAZlYjNWqZ7iIxJ4J7AVHyZwS2/9rCKResVTucDWV0DwOqBdIKna8YDnZstrXb19vmqfAAVhbwh
jjQ7Qf4=
`protect end_protected
