��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X���_B�v}|��{�� ��S;����%vtX��sf�����n|����XIN���>[�����_�p��̸��Ү?ո���ȃ6C˕ӕ���wl��k5���w��g�� b2	�+>_��l��w�4Q% �������d��*#��i�f/�N��&�a	���9j���	bD��<��_w��.��U����v�T\MV/�s�D����ZO��>9�	^���"������H
Q�n5�����7.R��)ќ�78�,��Ոi	'�#,���<z���fS֥i�	��oM�r�[���&��0�����C��m G��fޚ2eIL��:`K4�Y��3a�V(�+��wg��?,���+t���ȥN؏�>E�.5���UiW��0��M��NB~����鸪����=��YǤ��x�����%��ky�ap�+�g�� ��>�ɽ](]c�,�]�j����Hv��/��q��D����AҹR
�,'��7��� &޶���l������Ѹ2z��+lɜ����2�"ٗVm� 0�����o��^e9$����VY�p$H�o/s�q{��<�:�Ҿ�	��3|��e$���(ַ��U����z%C�@�k+��W~>_fM�Wj̆'3r�I#�T��b�|M�%~"}s�j.Q����,wȪ��~�}�P���y�Z���8�OҖ�gq/
���u�Q��܋�ׄ h��C�zB$yl�n��e���[Q��,��y:�v3M�<0vI#�Q������d1CS[3/E�F���T����tҠ�[N9^eh����D�#�`�@E��ړ��*9I�:_�8�׸��P�.l{o�h�oY�񳈬I���e.S���LQs�H|��T���"�����D�.}
�+0]GY�RPNF<�A��M�'��p3��*��)��ґA@s���l�3=�|h�}�iJ�K�ɐv��\�i��&�'y��9{{{]�ٲ�nI��~�-���G��;7>">�7����c/�;p~C��F� )DY�݉��"{�Ġ�DM�S?P B2`�S�bM���l�fw����V�Y�c s�+��-�C��Q��0dl�oQ}l�B"�o�Z��+ٓ�s�X�'����*.;pk6�&�hà�r��0�	��p�F�� �t��WϹ��ђl��E0�,��(�{~�Yx��o/2X��*��*�w�>��6E�i@]�!4�i^�ʨ�n��+�@4�z8�L�>�C'R�8=�c���8�K��\s��W~E��'k��i"���h�0��gZHg�;���@��j?�c�p�Wҏ��OY�x�Ȁk0��8������2�����+�x�g�~���gfq
,�@�F�	�b1��z���8@C���aτ��8O��:��Ԃ"ǭ:n)W΄��U�� ~���Z٬aU�"�NY��#[U�S�ϩz��ew\_d�U�Ѱ煴��/,?
 UT�-(a���V�><�8�y��̦_R�
Vrpx�i�u��p�_ն��-C�0��3�֟��P�0|�  -HG��zΫQ.&����D�*ֹ�"�»n%�#3<�ɏ�Z��=N��䆵@�,rc��$Z���xm;�J�UZMa�#0}Y�]�O�!}a�l����q<�Np2����ja��齓��T�O~��"OOK JN�ڣ��t���Lp=����'��9�Q��({.��f3���������kk�����%Z�5��~!�N��x>�%ye=<�}y�/>bN�P^��W\lȽ0�JAl�E���ē�hu��y��E�3���͌�x��6ʧS�]'k<�Ĳ�H�)-(�W�T.�]d�67��H��j�I좂���Q���pHg��'�ߢv��o�6`#�Ƶ���V�ɸ�<����r�x�ga�%�#H;G��"*�$-Sj?=gÂ���$�&r8�R#<���G��1a�r�T�>+�B����Hva�I��}���B7Y�8oI�r�ն����Z�u�a�F��5_"�D�M��D<Cy�$��s?�4��A l�e��Fh*��1����ծnO,mIz�� �M�V�0��)��G�qt	�I��4p):�7e���"�L���?�	e[��|Y�ן��G��6�R�z�Xn�Q+\p��;y՜���M�V_��u��H���t:��h���p�-95�t/��L�J,�Q����l�"=OU~������k�\e���,���xZ��~h�Y���=�rD���:�K��w���p���Ü�k�[ْW�b,P��VJo�E�>*��)5�T�L���nhDV����;L�&���[�,�'�YOSUY�^�)S�?�k
�y���ҏ��1Q5^�F胨��+\W{�%��2��zm�mn���Yv~�i2;;�p#�0��r��,�y�+! )zWF�������g'9Ղo�Èw�x�Ë]:l�E��r�p��e0���s��nOAѰfb��t��#�P|o	���?.�I^�D�Rs�~�Z��-��2I��gH��1'�/��l����G���p=渜��ׁpK�ۗ���ϓ�s\$�3��g�|>�c5��l�*	+��Q��ː�e��n%R�r'�c�"Բ��/�����hg��]�A�i�y�Rbb�,5yG���i��=��6��b��Vzf�r<Q񴤨�k}��\bN�c`�ז�Ț�g��ge��/l@uF�ƅ,N�T���W��Oå\k�����9��K����b10۫�_��`���o(���D�@I�� ׄ�g��[�U��q�C�V]9��g �#2[ލZO(Bɕ�fyw�t�^9\��2��
$�#pn�0�J�E����(��ꋄ+"K �{�Z�>�0�S �a�,��Z�N�%{��86�5s^kh{ʪ������W5�#+��L�<��jB�6ܽ���'~r����̊������	���� ��������g8��z�� �]������(���g��zjm� �)j@
W����7h�
��S�p���=?�,�V	χ0��p,���:��W� (C���y#-�:�a��Ս$�1��ڑmx����{��2Zsf����yI��c>QlL�z�藧]q���b&�ݺ��BO�I!�ٞw2�an]�g�V	�츘�iH�f�Ӯ~�1W~�7Ҥ��=�&��%�%j+ro��NO��AM��)u=��k[��A-��i�K�a��7.pp���@xQ��d�.�Z���D@�vz��u��K��&K��0�'MT�I��6�Bk>W���K��C�ŗ�
�������.ar���b��V.�W�7�i�5Pz+EAΠ�`5Pm�ag92�̩3c��S��b�>�d�|��.����"�"*�T�F�#	�W��)��	��m�j��V��*���>j�����衹k֭�28�649z8%��a��x����!J1��
n��J]Y�Pd�E����*w��}Tlq�����G�zl#6�����4�gj";=3�E-��Su����lI����[/�4ẹ|D]��i�B�[�k��.�jo^�=��'C/�P(��Ʋ��IgS���O ĭh�)���_/_��l�0�+�l��������˼B�䖐Jå-B}em�>e�Ѡ��rK��y��2KV=<�ߚ����������;'\H������b�����E	F����#���:ϭ�v��>�RH�'����pZ�x^�+�+_��,���6��"moR�`'g���5tr;",��"�&mO}�2 �0��R�#;�P��*W�f��i�*��Q-�y^�J=��w�fYā�h�	]�w�~\ �-����C���)̓��X����6��d�����v�@�{�z\��,��l�|pF����x&^���XY'�!8��&v��r�H�<PΒnm�L�0'��|Ȉ@$D��˰Ԫ��u�H�78��C��s�5�����ě��,�O��%��Kt��1������?����Ɔ$P>��U��j��l�)�!V��ϵ-zB�Um�\��P���y՘x#��3��ĵIXr�7'��%��}��|sr�wB���$�g����e�Q"���,@ӉW���l���H�o��K�\N`	#2�#x�սS����V`���䉅{���Il��5�2j>�s�e`��Yi*H}�@ƕ`�mU#�b������Ι/�Z�֬6��|�[���a{駿�ˮ١���$�zV�҈؇���+ "�0�%��
��qNcSۉ��3dq[w(�U��QDcN���8���~�I�n�W�6�Mj8(NI���#����A�Ϙ������*r��_�M��xQp��ir>⊤��&N�vn���u�փ@��T�,K(]M�-��']%-�(�����K>]Twi,�e\�͚���_+sЛ��Z!�v�$e?�n=���P��׊$��mj�����4��}7&I7�;��|v����}0;�R�*�B���O���1(|pIf�D�Y3��`�C	<6�;Ԋ"��K���.���dn��B��9>����`DC�#�rKC�~�{��t�kO(���~,?N�RC
��Pg#��Gݝ�c��$g�:���'9���퇾a}8�
4ރ���J��Σ����4���ELI����G�i1FĸE\N���ipZ�������<�����1�m�H�0���.��{A����'|�O�f����!�Uk��S��2ԥ ��R#����Ӌ���2����RO�4 �Z1PSJ3|�T6�Lდ���V���۹<��1s�F\�jf���H"$U�>�h����Οo,�ǩ��+���?�l���1�����]�'nf?��A[���L��Q������d]���K�����!A$ef����E)c���+�,�����#����������VU࿭��;!=',�z��{�~�1��IB,*9������XZ�����T(a
�w�"*����9� D���]�T�ؾ�
ƍ�Ky� {������N�����B�s��K\n���r�AtsE3�H �s�`��	��݈��r0sqڽ��� o�W'��D���$t�������^�@8o	GF㋆�N�j�r�(I$��� ���4��C.��CH}�Vhp�"��!+�~ .���	+�<�������Kg�W����窈&/����u��ə)�>R]����z�!g��L��n�[r)��|O^SΦ�Ԁ~�, @�Bn�Mr�9�2"J7�����W����l��ò�����T:��x�Ɔ��yЉ�Z�wQ:޸��{�n��l�S��Ŧ�9�L���n����GF�Vj�g/)��|�6�Y+��v���� S*Ozjɯ_����VW�P���U[��x{i����<�w�}�2�q�t�	%x�d��&6����
*�j�g�T�; �#�r9��됅�SjOXkbZfS�|�M�++�R�"�t4�z;nt�����[x�
5#�Q�����Ӽ������T��^p�l�[V�Z�Z�H�ż��-)�_C3}�
�/�r�i�/X�
�Q��Z�!L�=�H0�tቄ���5�	�}I�c\S��sǄ��:�H!�&�T�ȩ��Sr�4`�h]M�x��/9f�F�O�۸N)}?Ӣ��#�R����fa��.o���@Π�q��A�pG)�0&����F�����,�9l���"ʁ[��$��^W:��)�����/�PHy�q�g�2M��s������dT�VU��,�bqߺ�KY�B���gG��hdDck��7M���e�H�eXZ(��3�!&2k3b���K���ojgя�>�s�� ���K�d��{P굚�fo$�*0�4��:�c؊�G�zN�T��-���W�`�����E��Ք��S�Lڿ����op���F}$J[�lK��Ҁ�B��{�f��|���ҳ^�2R��tbH�+ǚX�9�]p�E,���h�֖��È�|u=�*ܴE���^���c�hzEA�mE�#aO4]���p4%FLL:��H�A_�T�v��Ζ(�!=[��c�K��hp
+�;PS6�:d�d����Q�_��f-�
����麣�8%�e������ur0ݐ�J>��Bݽ~�Y���4�b���v���E<��܆�/r�X.цY�V^RJ���c����X�����kb�� ����L��P�"�e�q_^�F�h�շ�^�S��Zү��DaaJ�u�ߓ�pw h�`�0/j��v��Yƺ��f���t��Ӗ�"^V:;��$*��sc����a�f��ƭ�G@ϻR:��εψ���FW�o�XL�c���<'�:�Q������qR�	���K*Tp�/�������^
*��F&r6/�~�!��ˏ���G��C�[$���R�����������G�/D���LT�K��U�X�����ۈ%�?[Vu}�H���Q����c��o��c�L/m�&�-���[���l׏�����V�}/j{�I� </�v��:���_t���T�Ė�=�u�H��Yv`e����3PfF��U|DpOߋηrh�����l����XS��:
|������^�S��È5+��q�)�����(c�Pſ�󿐀"�<TI�����(�i�KK�+��w�ł��Q]�w����N[8��@\�-Yot�Ӿ��UXȲĎ��`�w���j����W�VvX�yJ���/�M�����=X֏,����x��?3/�����[m`����r��m�h@�m��iz<Tt���͑�k���RBpF�]��=��C�і�A�䞠.r�/ߣp�*X���l�����K�X"�*�L0;|;�$�ک�'��޿*sL�O��i�f����!�-�`O�I�6�MW|��J�L�c	da�$���*����ଝ$4�Cn�R�~���q�C �J�GW�X>~ĬJH�2Y3;OY��;�M��a2�c}�1ZĪA��;	��F��N^�_C���Bb��h Hj$��~bF���#������i5=�5Q�PJ�6)�=�4��`�<�8�;�@���D{�}��U�G)n?����E�@A�#L%.ȵUi��)�5�s���Bӈ�!�ky=U
e6Us$�Zv�dA�����
ᓇ����o/����Ɛ��b�f?�#8GgY�V���\~��A��|� <�A�S>$8L�W#��XԑR���R��P̾�X�hE�g����<K���1����CmP��QԄ%Wyh�Ru/3�@���w�k���޾�$��8�8�u��^��V6P8�ĥU_"ܘ(MUN�8�ڳ������]P9�ځ!��xk�J���/�+�):Նt!��K���wF�P"���3��}]�~���C҆R�D\Z6��Ĕ�&�1�S�b�SФ�b��Y�>ݳᦤ�C�9I��!���^p�K���x��f(v��J�mv�H�]$=;�X�B8 �(G�b�m �^Z%�����߉T{��Y��⃁�&h��FB��Q`^;A`�Fz0j�;Z�5J՗�n��t:e6�	ϳ��oY�\.g�C���. voE�0����ױ��t�U�,�{���B4�z�J������n���o��W�¯#v����,��J��=�����e]\���S'J��Lv	B�u�6�����pű�r?�&�x���2��.˹
0)7���6��2�W���g�C��Q���k�� v�R`�0P�Q�	G�e{���d
⌨�X3��H�,���QS�!�����0e���%�+�e��:tJ��h����HhI���2��"��N��^I{�f�E�h�G��Y����L硪̋ꖽ�c�<]4��x��kD���2�.��Q���Y�ߞQ���~��~F�$g�-��У��B 2V]�5�����%S����t�2	U��`D�S�TU:q�F"ru�'�;��RЭ���UY}2N �/4R��|�^��R���;w�kPL!;��P�t�°��Dy9m?3��V�S�V�5"-X��3?H��w�>hդ�=̃�~3_��q�QJ*��\�`N�Zz.�*�4�{*_/��=�s'�Y�Ϛ-���d�+~	���T�Y��wկ�N̵@ :����ҙ�8�cӅ��]��Jz���$�Z�2i�D1�"+�7�f��yW��8W3{��G�d����P�HI�������j�6�9^��?�����=Y�l�$˞����h�Mz��\(�P=u�����gT�u�OD�̽��}\�K@�S�ë8����cn�R����N��(�"��$�A1�G:���O�%CNw��.�A���g�����;7����g��&
3X�1�:����jO�f@�	|��C���GOc�S���Z><��qc����g/�����z�=���~�'% DYp�-3=x���D�b���X�� !N�����#�1�Z�2�5>]�e��6l�����)�������xM���r�O!e95U�g���[4�V��L���/^�����E��9�����Re��ڡ@�̷~���Ĥ�oj��%�����2�8�8NF�*��"ǡoWR�w�d�7��%x����)�n�6zf��w���3�g�K����~�*>�h�*
���Q�}bS��9�C���NێS"��.fo^��
��(��]�x�������G�	:���L�Vs�.��
ڃ캧��S�?�f� X/�B��'�k�_QF��t8ppRH_��_h��k��P��v&��,�Z���}�=�4�ĕp�JŢS�7�^�H��¬ 7Mwp=�CukZ��V�w�
j�T9)r��Y�~���'Ҡ��y���D!`wb�9ܔ�����&p�b�`����@��!��Z�l�xE��2n�mn����d��"Mk9<�Ǣ�~�ʉ?���/��C��B�Y���AWeN�;�W,7��ְ�C�J�7 E��٤P�&B��n����{ �o�|�_J�+��ɵ��C���TSP��X��ܞ�u�~�1olk̶P�/b�5��}���:<:ӐZxa^�}"3�����E�Z����3�~
t<��UZl����r_ԙ9V)���XoK"��R�K�E#���kE���+��&u�T8���x3�=���f���t���6��<��X#j8�&�m74����k�p��Շ0��*��X��[L��DY��j\V�
����X4�+�v�YA�vt���D��X�荴��
)�ҘpoI��H#�,T���>?߿0`y��d6�3V������-֏4�s���9-(D��|��Z k���@u|������z�cX�\{kIc���H/�ټ�������|�������c��%Wx�2vd���+N��ԭ�D ���Z�G�d�Gm���C�`����n���/hCm��m�E�6:�v~�؁v;��:��D��>�JCA�4���T���;N��9�����jpnSq���0�̝_ZϬ�fJu �r��m��mA��)�x6� o7J�[�NՏ��z���.D���E��q��B�Y���Ґ��NI2�w����,�Jm�٥�[��,��	���5o����r҃�K@\I�	�v������	K(U��ړ&��u��|R��:��پ\�Y��K�:�&���Gq�	�aVx��M�\����ff�����Y�;���E$��بx擩�=�.T�fv`����6	<�rIA���|:��&�xM嘭�ל-��xk�ӆ� ${�n���OEPn�ou����&$� <��.�v���x�a|��F�7~?��dt�E�;���%�Jp���X�W	�@m4���<�31���1�%�I#d��ٯ�ː�O��4� �>�˾�@�������z[Irb�M���H	:�x��$�k=��2�o#�̹��V��3�k0?;ý�n��9�cB�+/׳9g�D�7Yad�7�l�9�S"ɅwQ�ą�v�9& VF n�lHa|g�=pI�s��8�r]�`�QE�hJ�@��� 6�����4��${����wxA�uX	�L��e$(Ʋ�����!�	������)���6 �p�61:�]��G��bb�@��2��`�.�(ո'ZE�X��6Qˣ�'R��rPD�J�X���(����˖�@1O����E��`��x�,��_�)�B�},�é���^�s�y���������m��a����Mݱ߮�a����U�<��˘r���s�L���L$ၽ��:��X��=�R�����i�L�p>POO]���_�`�B���+�a��xH�~�-@pȹG ����]N%��O1�LBR����[�#�O��W66M���=���������Cؒ:b����O|E�m�y,5ީ���:y�ُ5�0�ks�w�R7G���1�6B�qQ�nb)�TŻ	ࠅ$�1+�1磏�C'#YW�=`�F�!Ë����\����>�t�B��/���
�<��-gRI�!Х�e�z��p |�p��W�ަɯ}��O&(�C���3����Jg�F��Rg)A�O��}�)�`�$~xl���<��@_ p�|X�6��S�?�6��ѢQ�c�����i�T�����D��4LJ�K��h�=���޷l�N���̿��3��������܎Y�̈́�F�%�$�6٨*�j�?��|̅�rʹ�L)2��[�Jg+v��0^������"�I���|���%6X����S��MZh
W��h\�-��<F�:�؅�FYϋ=j %U~�+_�:����7��ش��embx�an�ck�!,b��=Ζ���+����)s Y%f�~�(�&xl+L���;��=[uPfZ!�mm�F�*�����H��N�C�{�k�D���GB�<=U��p �V��c�[�H~�;lnJ�apO��*��{/������^mց��na�h��[^�)�����GiА����8}�8�i�}���j�hl\@`ό����2���J�vH���]�Mm`��JZ<��o�(���߄�=4Q�L�t�'��/2�>�����9��b��(�wX�`V���͓ �Ұ��5��wQ+�L.b���T�+%��^8N�%f�b��9��"�h�{`���'�,9���~F>��T�84��y?��3��������)���n���@��,�i�o�(U>�]����r��B�Q�]��}.k��}:��z��{F;U���96H�Y�����[��ɏ����Q�������D%,������z匛D�ʓ���r�C��t���L���c$Ч��]@.
��R��_��h서��2��׭��>����6�U���mH������yic���ק<��~_܁O�+�v��f�(�X�����mS��/�����2�jn6���x�E�n�E�J�x:wa�Y?�ݡ�$��2tcL����Y��"j�b��P���{� ��D�f^['K�N%��3hKB?�(~Y�ykܾ��%q	�N�1�/~�Tylr��#�x�q��7.����ְ�2���ƭ�B�1�� ϱ�GT��*��(2aH�r���&�P2�_��B�5O��#��z��	Q���
�x¾�RJvI;	�cc�Q��7Y�[cߖT���:#�t�lb�	�Pv
�Ŝ���6��Ou��{P����(��a0_�����;(\g�1KT&l�*"�����sͰZ�"iǿj�1�.u�*V�-0�Q3��uh�X�ؔ,�
���Z�G�X��Y�W=<�7�h�����F�j�����+q����� �m}��>�@ϢC낫��k �U�-�g��c/by3@V?��A6����gSiq�#0,�#��D��y&��{5O���<%����5�(��R�m�Z��/7���csmI��\�p�MA&5i��Xa�7xaGR����N���Z�C]��lGx!�.=L*���SB���Xld���4h������bt���7���z_l��K� 4�y4������y�+ U�R�`P�����9��(Ĕ�LIɵDЇ�߁��HC�8�����Z`��T?����JQ+讌+2���w�r���=�o�� ��֫�V�Wv�v�%ȞD�g���Pb(��wl	�������f���̖D�v�l�#[�b�D? ��\[����#%}�a
R�S�;�?7X\�SqR���m(y��A2t���!�qJ�.g{��{� ��d���+�����o2lƯD��ߠ6�,ڔ�Vs�����4G��\H�����M�GPM���4a�Q����:�,��SHi�%��S��RC�ڠ>��>p�)�,O��_��:�#j���i�k�k>��Ƣ{ý��a�VKVL>)$Ȼ�"`��Ώ]�7�PG��Y0�42.�_p1t%�GPP/@cpy�)�Apr_��E�=����`�~2^HfB6g��C�32v�_[�n�i0��%d���~�z�����<�\]����0L�&������Cm9>#��]Ю�F\/��O�Ћ=�X� o4R���-�|�^�y�N��M#��4ґ=ךX"�n���y����p�(�j��/a[������$!� ͼ�JU�F�Z�{�-�t�J����K�i�΋�v6'���W�]r#��H�s��O�D���p*>���Hqh@

c#��s� �3�t���zZ`�5xL����i���ׂe�\jH�=�WN�zu�L��;C�e��Y�����=�/WX���|d����;���T8���~�N��Lw�89�*��;	� =|@'�ϻ���+(��j��J��?/:�ע#��0�HJ��Q=4˂�]�t6!G��i���T*�~\N��#�#�� q��Ө����R�Za�g��sC��ZL<�c
L1k��C��������>@G������5�s�,�ՙ\����/2=��Q�_ۭ}�S�}��1 >��,�K�ԋ�S���8j��%۱;�l�דx��$=y�!ΧsL��g��!�dV���M��[1\?��������`�Z��}mj�Gȩ�"�~�Kr��h>N�A��n�.��xv�c`  \�i�}q��~عEO-{c��w ������ԛ�vZ"V3���OU��8dOxG�*<���mҮь��P���v��4?����F�67S�D�Y=;�j�3B��?dؓ'���M����%�.0}�]�]%MAOɟ�:��=.�5%��t��yjU)�̗��Qj0���Q��/ХFYO[��L�a�QA%G����n�V0��q��0 �Q�Z�L �%X���b�
��jz��}��I���9<.��rD,t;�����#H����l?�����	o�\�`��KH��g���($�!��\Q2�	H�c��J�e��-_�\�ct��-z��o5\#��΍���3r�P�X)ٙ���WY
�sm����Iu�fV�g�DNO���/8Z��ۘ���P ��}��\��J8V�R��H�՜ن�@Ŀ�^������V
��Pn"A j2!G�0��@R0���}�O��Yv˓��L&��C���)��[��ku���eY'�7�ٛ�+�i��2���0j�S)!�Q�1v>����� �&O� >F����%j�E�8uұo������,���[�I��.I��_q"�চQ�	�q�J7��Zۑ�lZ����+I1��m#і��CU�Q8��\tCjysN�{P�sT@Q����BN�3k�u�`��LH�3پ���9�X�-����A��x�|Z�)e���:��.��Qȹ8�눮�����rC�حg��V ���yP�1�^}��=�z|7'�D^`e�,h��O�Pf��|�L7���Ѹ��@�@��������&T��ő�t{p[���:	�;��+��ym�t��݈��w�Ae�$��O�w������栅5�����t�ط��.\ �ړ�^�E�Zߔ�b70\�"��t��0޽��W�6��~R9�p�F�n�\��&�om��!�[ٱ`ּ(L_���lC��������4ٲ����8�T�#@�=���v�#�jlH���Y��t�	WbM�l���d��
\�a�����i�;��Oٖ2 T��|����ĵ��z"��/0&�-I�p�a�%�7�6��8���0V0f����\;��M����?l&���R��G�lˌ�)'��u6���g�۱��f΋1An����q�gVOv��q%D6�5�ؒ�h�r��S����]n~�y���C]�����HP�s�S���m���������d X��T���]����>!��s��؄Y��+�����i���MZPkZ�t
T��>fӸ0����˽�h���.k�^"�l�$E�|N��}_�7w;��ǞP�w!@��l�J$T�����H�},~W{� ���=ɏ�}�nq�wNb`?6��ԚB��YK�p��P+Oދ0�����ڍy(�����s�Q�e���
X���_�9$'o������3\�[̟h���3����G���*T�-�� ������Б��+8�5��^����xN+��<i��{it�i���r��
!�[�ܴ�fe@zUD�&F`���܌�Хcc�]���h�V8hV:wA��;y�밥72����]j�bT�wq��5p3����1y^�y ;L���i��72��-�Z�N~7�چ'���[��c�������$�D��@�R���D[��}n٣Q�����+���jfE�m�9)���JAJ �Y/4_�h�PG������(Z�4���Y�4�Q�jM��� !���]�|R;ʒO��B���/*�Ym�zdSU!=���O����83�=�<AbӦ��.�#m�Qb@�k���Ӿ�-6ΧnvI9���	�`_�4�D�EVy��#-�
�jOP��$6�h�N�FJ:���OM\h����/�C���}`LX���'�������U���~h=�ś��I�wxF��?�`MZ��+�����(�������*�j������ �����vT����.a�wD�Oў�v\�d^p�����o���}�(s�|���B�B�ȗ��������.�5�,���n�} Ԯ�%�@_4�N=��#<m�����~P��U �F�`yScu�~���������J���`m}�C2י�R�A��L���g���fs�N�����B%�)k7�|D`�Ch���>#�a����w�(�%1ͷ�ta�@\��W���]=�up����.o%7t��o����Ŷ�j�c�EW��p8�7t��e/����S�i��Nd	߫��¶3�)�S����nx�!��(�Sk�{bK�柭g�ـy�"R�n�}ed���Z��a��T�IF]i���r��K�p�Md�ۧ�ɶI��8��e�΁��<
��\����g5�T������O�Gx)�O�J���������|�`6�P�[��W�4kD����<�K z+]x"����˃����;�'a)���涰8K<?���I��mGY��C�f	&���.�oai,
����k$֋����K�����ş���V�i�� -p�ѳ5Ƶ½�\�j��A�u,~@���Ɓ�֦19�i��1<lPh�A*�M@�:qv
�W}}�x�pջʊP�WX�`I�C�%K�p��Q��@�z�<�r�I\�h-���: ���C#F��d�F;s�)7(.	�W�u�6�>�K<pa����W9��E��CZ��R�(�kH�㞐)��tٓ����m;<�b���#�t h�A(��7,�؞YDױ�"��tJ�r5!s6��G5ه�*��������R,?�:���Y�=�L�o�����Gߜ�J�T m��*��zt���2\F��W�ˑ3�Èh4�g�ڔ3���-W���_k��3�6���o~�Z���g�`tEB�?���5�D�1c�
(Ji5��%n�ɒ�m��z�bͧ n�~�s�.4e�9��&ˣ_@�gEo�S+���f,'�M�|;� qS�dܷ~�����B��x�O5�*T�=B<`ͪ�x�FI�-֍�U�zj�<�[Zym�G^��Zէv�	�D�bN4��g��".�zb�E٨��	��Q�3W[b�4>Z����ʶ�ʯ���m��&�-�����Llg���~i�4�$R�Zq�͝I+Yg���r�0�E]ݲ���[�2�O���u�X!?��l&�2'�W���߄���-d[WK1h\Jʖ�e�3��ۃQm����V�b�`u�V�4��|��	�9�l����� Xǒ�r[:�ٯ����?��.��%���J���'�8�]���-N.�z�H��H¶V
�9T�Rҙ����ϫ=�u�l���7�L �ST眄y&î��bL��:44���Aۮ�>�c��׏�6�a]�m��ӝ�wp��}B�`����lmo���Afq����c���G0p#��hi���݁���4;�Yĺk�����5{�`�za�N�� _*�:�2;��L�Y $8|	d3��.���H�������;�8}[���fw����Vk����Hf%�i��$D���3 ��,aY��)�Qc��TΡ�݆`���3���E�E~��Ro�"ؼ�ۺU�N>Z��>_%�i�����o�,�b�,��	�X����/�T���JZsA�$H4�T����+5�E�}��B�W9	R�5�J��l�D2������q}��f'�B�
/1P4���*W��&=�w_�Z��^�6�͐��{W"�SO˩�B7���}5!��-A��Lz�DLVA]�����1��0([˾����Y��GY1}���.9C���}Z�֭�v֭�F(�\�~�0i���ǚ��kmR�8�����>�YD��v���֍��ִ�3�d׊���P~!DkL�0<pz�H�z�l�����k4�ǢUU�g�=��5Ĵ�__Ʒ���x����޹����>�5VFHJN�N��]O5�)�����s���8�~NKf�4�]�K�"-j!�+,�:E�O&2����"$5���b���[}���X��f��c�-���1 �{'��Ty��F����լk�;��V�x�/ �!�5I^)Jr@�p+�������A��$�"�q����7����&��}I�l��Q����i���_�C�Vu7@��,�}���Tc���r�j��_H<�#I[�sl�u�0n~#ۂ�)L�a#������&&-���������	ՏQ���_�?s��w'�ǥ̹�'��|Q`
[�Rԕ�b����c��+�Y��N:��#\��>5$r�Q��cP�h��m�?��SMߔ{4��Hk���e��M��Gi�Uo���f9>z=�][E�^'8��"}�O�}>tU�ϓZi!�$���❛uz�k�퉢��s����Wh���,�~�kNe}�D�����4�>"]q�������ב~=�)�oEkh��@�T����pD��f�(�F���G5��x��ʦ����!��Zt n�6������U� @�J-"�t�oM�!<�Ҵ��ϰ�p�O皇�`%#{zVY�m)7�y�(5��=I��A���{�w� W�[H̤YQ��7���m�b�V*B�c4�Օ�1��ͼ\3�L�%�t�өݒ�V;�o�O��纪�}���_~��$��3�2�iM�9����'�ĚS=5s�-�eUڅ�N�b��۰_F�U�ܹ T������������Ez�M�}9k�����G�}4�Lٍ�=
Ym������~~Y̔7y,S�� {^lhy��́�I����yH�?�4�L�D1
��h_�Z���	%_��ڌg�@�c���.��Cw���a�%���cQ���ސ��鳝��A3��Wo�𑡏��&d�j+�,����o3j�6��]��Oc#c��|M��y�?�M�ub Q ����#}&�O��
;�zf�o��H1"I����N�bd��Q(xSxF����.��{,0mUk�1W�p4s������c�Vj��eP���хz���{��8�Z��o�H;ͦD��C��>�jY�Pn\�dn
(����d}��חY�Е�J~�/��Ё��ܮ�"~h�����I6��E��z�ࢎ��P�@C<��De9���B�/�_��_M�̵ԩ�C�C_"_\���A�7�{����ސ���5(�%[A�8I��\�9��3�ԭ��}�$�mҵ����KH��90���SEZ􉬣��D��]z����(�`Τc�M��1���3����q���w����� c$�4�0x������p�3q�g��y9ß0�;mf�����,�a��6���[���`�5��R8�6�g�Iv��lۖ�a��Z�N=�	O��-����`Nc�A]A~g_��"d����i�T�P$B�b�1�>e����p��l�0��G�y@]/�z;���5m����{޾��I*��,8��q��Xҍ�R��w,�W�P.�A|n���i*���E~��^دt���������Ap��Qx?�-9���=:�q��Q��{���jLz�iDO�!"�`2H��ȧ��q�����*
�3�m��g��0-�c���Go�������ʆ持�����v��Щ����G�B�z��X7�[/S�Ɛ\��9�E$ZX-Q/V�ɰf��t�H��?Hzs�:��(�j>�U���f�����)J�~m��m�yQ�V���2}<�'L1A'?��I�pW/�� c����9��\�u��= θe��Y���v���t�
��JEx��L����ƲA_�X-g�6���C�U��@[u>��̬���e��]����Ǌ��h����E��L_����Š����1��:�W�Y^��5Lh���\�U��x_��EP:��v9�%
~g�R����O&'��m�1���Y� s$�bN�ܽ�:�g^R�4?2	.�3��[rn�V	*���~yE����Kh�e�]��t�<ϯ0��d*�|;<���#s�E�C1����f���xe�'�T��H�e�YC�)�Exx�X,c�.��3+��h$Z�}�cvzK�`+k�CQ_͏���z�<K!�l�U"`a8�`�U �Z���zo��î.
�8�NSk��يN���� �ͳpx��8����O/�ueTV]�t�?���ƛ� ��?CP��r�@�l����ۼ�� J��+E�T�I!^�9��Z����C+� A���9h��ā{��B��*�ѻ�QҤF��4���`k�N�!ef�/�C-_9
��|Уͽ�X�箪XZ�_m�֋��]h��!!���ԥC<�?�VqQ='��F�Q4�,x<
]��Pۍb"�Ogk5�s�O��9υ���i�n�!�v������&�ez�px�UR�W������:�H����BsO:�'%,��Յ��C�� �����~H�n	#sI���z�԰GPcxˋ]��_E�"��|�H��l��Y 'w6�X��,g����V��B��1��Wԧ��ZJN((�k�&�{�vG��êg~ �X>�X�6H���Q�TK?���.��[+�4N���U�(d�LUb<h7$X���c�,i.��E��죬�� �!��R�f*w��J�TJt��k,c�_��\%b|ߌ����#���O2����d���UR,\`[�V����<��ú��OM"@B�MД�8|Z�U�K9���0���]b��qQ���ûwم���\�Z��e݇(���L���s�x*1T4�=E�}m���k��"�"S��Ugaa���u�&��6����ߔ�^��-.����Qz���z�-�meft㯬�r\�n�Y�̽�StR�>Ic�e�s���/]��L:������p"H��sD�z%�$f�+(au��K�����J9tiLqM��+��-m�R��(�5�m��B���S˹�L��4(�vw���҃ğ�c��S'JUaA�|&��G�Y����������� ����/{��W5�0����z��9��0jAv��6O�
f�v/jchi�6(`EA�[��qG�|	FJ�v���Ix�%����uz,?��Q��D.'j꠰�C��Q���-��|�HdV�����Q�����L�*v3����o����^nw|1�әmk��z۽�D_I���=���X�/@�3&�gDD�����N���}M��w��2d
��X��R��ĩ �pbp]��� eE���^�s)��8�X�;Ù����{�@`B.��h�/rͰB��j�R�ɉ������ɇ{��D����-�������9�-��jcG���*�����#z$�<�EB*{�����	B�F�F��Xa?h@���A('q\D�k$�W�6Q%E��-��Z��Zs(��{��~�#@��YT�����)ke�U�%�G|�-�N�r�Br�!9�za\��O���Ơ�Z�����FBJ
�G���`�t�X�+�on �zM��Ŷ����i�������w�y��S�)|��.����������_����v��:Hw�`[�+���ܟ���]r))~��A���εk'_!כ�$Q]�����(��c������(K>��oQ�^h\`�@�?�eZX1y�0'���i9A��Z�e��6ocvZ��~���c�Ӂ¦�����5QV �*1}xy�˪u}�̀L��l�!`O��;�r9h{��!kA>�����3��J"&����[���X���Z0��̶E�F���PT?顉��pؙ�Vv�6�+)M�����*����.\��C/�m�m:H��H0��R.0�j�����#�� tL��O(E�8�a&��Ӣ)���ȑ��&	� MY��3ğ'ή�_b��>�OB�q�<�R(JjӹE����W��/����F����s|q'	��}��on|yt7Gh~Ӈ�!�I69��/��q���W�����H'ca�:����⓺���� 
������]��p`�}�_=����R=�+����9wq�4aƚ �X�d���������"W���`~���w1
� "Q��<Q���ew+%�R	�T�i��>�Xk����3"gm���d#���i�X&o<YX�	���� W�J��W�������e���U�2ى�޵�Y�������=�,6��V6b��T�6����	�q&t�,>e0@#�߇�'�~a�������[�#����f�~�1��S�2��6�Y��i���0��R��2zW�1���z�F�ɲ�Nk����|��p�$,� .?M����E@���'��Z"Ha�
�"�����\����t×ƴ�:! ,{�g��د` �0c�=��}�:����;��x���˖Z��8�k�M����O6	�h�ET�ŕ����<[��;u���^tj�����f�و�]VݣiK��M��=\�]qd�ʪ�+�h{�[Rb�Qv�),sU䥶O�Ԩ3�G:f*����!���B�����'''�쓱��! v��M*�Ş5���!�	}�+m} E����"����J*�4۹;҇�Y�u`b�ye�Q��f�i�l��[ۢ6	`�rib��� �sf���q��	z�"�ɍ��*�G���=�x���>L�%'m����G�ϧ��Ғu�,Jev���?��o� r�$�Y�ߣ��>���l�l�*G|��M�9yuf�+-��d��S�PV��J8���r�Ѷ�X6��:�Kr�"&���$�&"9{���4n�P2���{6���u�G�~遐����vA�����E����ݥPGN>�Y]��&:I�|q��OE�4іP�S���\�' v��ӝ"	�5�K�y�!���hUw����s[CƄ�4�0t{�T��b%�8̉�`�S��KqRk�̢�j<�3�'p}��F�'6�� /�p���gI�/�Z��&q�ƈ���{<��1�%N��k�R��9�zOD�����;+[֫6ʞnv��i�wy���ga��.2�� �\�H�?�$�D
S��D�N�7���N^O��;��jQb��.�!�Ca&�?YG3�	�ԁ㏞ R)�Nz	����{ſ|o�k���w�=D���"�M�5e��zw�S���P-��"4�O�kϾQZ>��nR^�C���^V���-&2N���#��+3ؤ��
�C�U{��3�7�U�ɃBo�?ݓ�V��;��,m��8�(F�{�c��Q9~���ApdH�a���Ξw�G09JGռ�PT��X>K�2��%�1�^���Iޘ�B�nv `�#�.��<���p�޹���u�)�0nk��p�KT�?m���]���jt2��U���W�<�ٌ
�8ҧ�nJ�v�>��E�_����)ң�l[��Y -���O/O�|$Z���Eo�b��c�J1�"�b��;r=��l�쩣��3�����:І��`��Ӊ���ú�$��Yd
p-�0qc�,6�C��Hը��+g���rG!P��{�h�	*H��e�BH%�J��N6!ݿ��y֩Џ%�̩����L�����̊~G�	ԭ�w��2ɤ��I��Oh11��{�T�b�8����I!R�A�����)).A�q�;�Zٱ�Z���J�r+��]Ej�3kd�ɔȎ	�IcC��sB�'h��짥`h <J�@��Y�9K�EI��J=a�Dʜ�H�(�D[Ǟ#�K������,srǯ�b�V�VX'��%&\ *���N����P։g�/_A]	?�KN��-Q���@đ 0�֣{[�����J�i7<�#��	njE��䉢q��v�Wd��Hx��[���.�b���n<Z&��ڕ�dM��>��6��V��~�f�N\
�ݍ?WD�'��f���+�����Bh׋8�j������GU�\6�#����A�-3�}Z�Mk.u٭ #%�ٽ��g9��_��.AŲ^x%d��2?0���&="���5Pr�m2��Ɨ\���%�^L�����^�����餲̔�\3�\�Y��vt����f��m٘�G1	>dY��ߗ[n ݕ�X�a��1��
�C�3#�ً������ǮQ��y����xT�7X��Ȏ{ۂ�s���HJ[H�1K��3��Z6R��;5{��
�������x�@��#'�ꄀ�7������=_�W������ʕ�Z[8��&6ҝ��Q����57%�< K][x}-[����_X_'�[�V�d�-ntv�� F"/�[�X�������k#gYu�]��[4��.�qҧ�I��6*W�Ӕ���n!"&���rŜ��)��3��S>�<`QL��=���:�0��'M�N�G��T���)Y�v�����iM��CB�;C@_[
��#�EӒU�d��S�/�#�F��rŎ���=�T��.�*�'���a"���C<����'��X�/�-��}b� I�v�`KI��$�W��d�����cw���ٛZ2[{��{��.���`ʙ�>��An"iY���������k�8��$A��K*�T�(�P��� )n�������LO}���n�O2�yl�!l�����P�[rkA�J�.��\ںE<��s8^�%�f��M��v��m���C�����E�'e�؜*�m��tSZ^�H������jN���/��O�#A����nU�����;즂s�S�#��1$N S*"����'[yMw`�7��uwm���aT$�xX��N9�}ML:c�%������g��1^��d'Yig(��//�f��,�ƇY��p_q�Q���F=s\x�&��a7K�[RA_�v�б8뉇���� ��ߠc��������k/�kK�A( �n=��]���������bi�H.i�4�q�K���5�����T/[��j�_W<�X�o��~��q��t����C�T�7Up��M��&[մ���H���2���ƅ�kP�Z8o��@NS���lh�i�K�Oϵ5��gtc[t���`V��5��g��P����qb{%X�"�nR��ά,=���w\����{8�}��$��e�#^|4��9WB���>����:��=�A�iN�A�����WǓ�u�ͦ��n�p-\	 ��h����Gr_�/ ���������F���������W�w3���H{U�J"��"���i}�E�ᧀx��t�o>.v��ol�X�U5�H42�?T�8�iZ��X�i�	{��?��"�'�s�? �O�1v�@ �ŕ+���X�� �1l�w�V�埢����SI	7�2��2r¸��.�Pi�&	�\��k��d������;�ᅷ'Pa�ƋI�h���?K�31�v�,I�y�Y�f����Ǉ����o5��UW
P�巂��d�(w�;��nvS��4l��؜~О��&�w��k��?H�U����
�U���I`RMc��r�Fz���U>�
���2�r�e^������%he���<���ׯ.��)�����<���#N«?�-��y�H�צ��?���51����<�L]�[/��
��(� ����V/VTT;b�|�|>�o��T�U���]`a�qw�lU��<m����J��K:��U49�+<��N�0�VϙKIy�%��S�m���:�X�R��lɖ�,�;s���.[�'�Kx��ӫ�B�U�Tn�'�<�O"&� ��G���w����H���2߄�{v�S?Kŵ����Q�^$K�S��|��ɿݨ븕�{3���fR�̐D���M0{;A$������ޅ"��!O��5:b�������دN�JQ��ZO�#;4��#b�
mN뤼�҆�3��u���!{}���~ʂ+޿ˠ̲�m7J�2
�SҬGX����:�v^*�\'4�M��+0M�l�HS�Z����,k���X�ɇh�%�m+��,J���a�α�_��u�&T����@��|���I;�J�^��������oi23���]*��|��?;��ȇ߂{�kb���(��&#|LqLΛw�=���#�����q����bz��0�%����o�lnUh�&��Y)�K�ʳ��7IM������ߡ�Z�6��-���8lP5���8�Ȉ?("�#󨅖�e8ǧRl ){��y�7f�y��S�B�g�ӵg�ۏժ�h�&0�YQ�h��V��0�����F��� P�mSW�͵��˦�5�;��t�
��p�n@b��4��?����7���פL���6����u���¢̣+�:���b+�~=��.��i'a��ٮ�U�"f�'�\��%��o�X���4b B$�<�0i�?�g�u,�:q����,vM6q�,����l���4L�Bk����$!���DK�W�������3_����k�..��6��N��`�e�CG���N#�km���c��ax�\J��o;=����q�f(���m>`BO�2�S��Y���r�+�[g��z�Rx�r<�oP�QA�G��#E�9Q�@��(i���D_@.�T��ž����x���X�s�&_�x  ��Z6����p�p�C�Y���yu�GbOZ�}�����dm�mW����"(m,h(~�
�d�0^��%��� h;R�#�x��4�!o�
ʱ�;(=�� 9���hJ���K�q��;��|�s�� ����_���HY�u�������G;Mtc�>!�26�'�$�4l���2PQ�!�U�}���B�vT�Q�> ��{GO�@��`J���L��aLE_9�]�iL���U�n?)<�	�2��y(�����S,���
�{yw[�'��sL>��	�?�;�װ�dzWe��*Q�سQO	ue`�l����EM����c?^e�~��I��ͷ; Pu���_�o��2�Ϧ�Q�n(%݋�FS��6�W��k�dR����x�9x�wo:f���� .}ux!0U��R��vԉ�����w��m%O/��hLE��(P�T�H:��P�MRR2z0G��m�����x���^x�j����-7�Iu;�g֛eB��(��St<;�E�kM�8l��� ��9�1�Y(8dU�����}E���!�{���������S}��xᲸ#�N�*O'�#�����Of�rpI{���E�%� -o��K,��!�����D/�8�o�Z� f�����Q�m5')l��DU.%ӣM�βs:�Ik:|a��'��H$r=���@P��K����۪w����������h��X�����>�ȍbO��Mb��?<#3=S�����+�o���b��vѓ��J�!������Nf��7�`���'?7�L@�J�h�r���0�b��N �!���4=q.����-�`� "�~#-a�z0�s0�{�/<�0�PMqW��n���G�Y#�Y���X
Z��:f��v��*�2�}m��8ޞʔn��L]s;jS�% ?��:���5{��V��dl�>ê\�k�V&����@�֘m�*e�\����gr��_����CtKN�`;����<_�%�3�`�c��j*������[�1�?�3�H��H����UiƁL��%�)��<1o�M�P|)�ğ�/O������=�[\�1��$WY2�SB�Q�Ā��xѯ�yy��!ڍ)�`Y��5Z��b>��Z