-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Rn0j6DRylnUjtZ62fYJjM0RflJenWwPntaOJWxOLNG9mfda2oRYeOfoFfiyCzFFW9JjYUFPTFbnq
plhMB9OovRjCtoY2m0sArXPopFxY5Vcd90Phf17eh4KThHxkTorKhIVeOlFTJaESQ89GMUobj5pA
z7rSeJFHLKnSvF06nq06sS9WMNs5qQJhNP0KZoScMlcu7BnoptSDgsW4P/jGaxSXRcCJ2TYpjeni
QHKz+d2v37umWnISkXvcvGQbB+DYIDIi1FmsD7RCe4tQC/IuUpvFupTwKIjNkaWWxIvzRQTf864t
2lmv5dP8I7gmVC9n/DH4NjQa5F7+IqV5C1lHYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
wAgygoHs4iRgiN3mKfOTTr5AnjmvSMOi+37pMrfkM3G8HHZUpAqoYXfRvwQ4AXuA48WRobl1wygm
szYZqYH57HMTrye+c4tTXe7SAec1k9rZcahPIUyKVx3uP+hykCqvhF3rZyROjdOHW0wutBjCn6zH
ixr0YdnK6gleRY3eUWGjmSPu/K3ZUUCZvzQCCy0222Z6Kne1nh0X2VUeewW6dH0BduAQ+BFc1qvf
3txVmcq3aLkYCdXxmgB/9pClw7aGpaTTaTIOgxUhf6R4VU36b2NwAY63y3olzIrG4XMu9VSYi26p
YSliVy23pD0PpxU/mrdTHoBfXIXKzn70JXuQFY/q5YZbZm1XHh9JITgFRH2qCWs2VnBQ0SfvB/kj
yW16LmYeLLlYnSfs8WqWBUua1oWukOZ7vBL76FmuJbXWqVkl5YpELXvEKBU9fYUDha75p94HhmVS
KWVLk4paAhANRt6sRMJyz4uLddCdmE1nrGM+zjEJT9X3Hnm34LjqbjQS09DwS61dK7QOvDMqe8nQ
/RVVPOquN1coeXYZMkfHmI3oxDJfQ+JRXXic8pgB/dKm1KKg0yvBp/Ifcu8tEGLyXjzjuk79hVfo
q8nCPC3yZhABs13hhejDne5J40UZC+4e+LZYjB8nzkNjvq3nUPXK5NB1+LrFaC54GbIEv9Gu4zs4
w4SNcTErFmMLyG2jnIQLGLhnQ9mf8EBeSRn+PBcnoMR5vOoEu9jVK5qqUw0TltjElC14wlK5WlhU
E+kQwwPwUASxeNWJkdclO3DPlQub4kHO4w0rntARJM8acQf8MO9vhPD5N37KoiL0lTNPzCmU529/
whBUoPkFRTYolsR61jOM+0aW3ElSYMPDjcefji/vo8bNFJEDw+1kElsgddAg0XKyv9/q1htnwZz7
UxxblM7up5aCV1D3nfOulkCk4TP04D2+USVmSPSZrEHVfpuoBVc+gzYZo6CdJKbTxF6Y7CqBezn3
hUHtKy3doR+lOQdmTId5g8cqeSt3vXngehDOWiHxKwsUqrojQGAv3j091pN+8P7IEYAdG6luEFpA
z0BCSvZNcvAo/uLdLl8eNJUtAVZfwX6JyNE3A/lcSGEIgao0pAM1BL2PcNpZVcg4cCnplsJVdUOw
vRMudqEPZqCBdwIRa2kBSsV+Ucn3WZp1CPGzvGFucGZCcKp/4bfvaQQROCjc49r9BgnAJIDwAY8y
jv2eUXCggP+Giv9zqYaYohsxSggEZBAsQHIJ9brf43emU3ohlsXUpg1KBj4JxI7ohxPl/nb2Rn1Y
w53DDwRT446ihFc6vJ8LOTkpBgBtm7sVjW/Jy9hzL4j+HdwbQqkSLA5WNJimtOZqLEbdFkzXNOgc
IBQkjoCu+VHRmHuKhWBe4hu57rZAZWat7ntRnfktWirEF+bxFX1+vLu7TgT4cGislYA6YNgoK/9d
PBr1OI8S6oX38tEOB41lIO4msOupa26XKzkuuPgiK6hQOukGt4+2uxvR2GMMyyAMvLsm/TB9IDae
YYEwW4Rd5S0UxqGATh/W+M0sbEVy1VVZ2Qo3/WC6MYt/2txd4TVe8kgJgMmwoc2taogSfnEgSYP6
PoLiPx7PVPKV71TJcnqcKgTYpGX1d/VMwLoIX2BDX4EJeyrlB+Ein7gSPdm5XbYzDplwagbU6tHd
MwUQi4V4RTBtKw1YmsNKTzSFRtzM4RAsVrqkU+D4HEWwaQ3P0TDDeLv2smuhWqLmmnI8eX8sjMPv
NhKyDJub1mzfnBwipfXjiuJa7gh+Bm+58KmPr6+6rro5F+11pZ0VggPQTA8cTCKICgdbabCI6DVj
QrFoXVLErfmE3tkiRPT2DrvWxmNtoAmKuCler+a8rjpHHfkUHdfnUpXmvDvlsWupkQjlgjZMb0zg
nlYD7Pjcl+4/kjymkUUqvH0CuMPZHencj7YlBb30NajQGyxsoS78Rj1r/yO18XJurgdT+apdJs/P
BOINnnqCNUz6VkYxSCLEVbpEy8IgQLQLPNRYJfRq34TdL9WtAgy7zvN2W92bOnPO3pTm7eAxBwZz
zJpDHaIlZLyZ0NyrDc6h7IzRaFgKA1w9UmVRXtObpVAvrWOxgjJZRt0IEOci5hVAGkykffrzZAlX
J9w/3GYqt63iRAsrblFFmX1dcpOz2AIeinBRcnLWAzTg3N+erM7vZhaIAjiIbvUEXqeEZPBg/ppZ
x2t0Xw5oOkn396yGrqZsL9qGg42e5x+aI55hcLRh5k5hGufZuw0sOgQE0nySq1Bn4ZjEZ/CwSd2K
p4iUOvcf5mYG0W0JYKyh1xVdv4VUM5TXmO/vZD+XLZ4hLzH31WJDvDp7LDxAD+09ozVX7F0T1OuX
FfT3R+B4OXfEja6HtSvgZlr2CFU5ckfE0YfhV8tbZ9uHjvsWPeJnXMFE78tT5u8PEE4NwKyTFDn+
BuV7ZoQwD7TwsWP8sRgwIhMmYCshwbfzdqNl2/E638yaOecjOfYpBl5Hh/WpuuIWDxO/IN+1u2MW
upXCE6gjz87nZGn/mfihBplulhJfqNPNlcytIuL8W1EVAYqNY/bQRhBmgdF4/QHxc/6D0vA6nilz
d9PukzbBzlBy9y8GpemXyg6gb4zihCdAlxZU0y7w5hzMqiPtkgHTG1+uK5NTtQpoLvKDTW8GSZda
3gNfu0EQksYwt8OD4UpsDgIm72SY8q8rleQ27RVhxHN8eO6lv7TP8i3C5HJlyS4h5pLHftICNq+p
LN9OC7JofV/C1egeoTGI8lDLUqDHd5gUAO+ND4iet1NGXntQGR1XX+m5q0kuD0ozCx8Rg/R3V3tS
7gKdCANYHIFAtOFC58Hz7VgOzox1PgI94KL/73DB2JOTbl3PI6p7BHkjCpNV75M5jKIv8nl+hX2U
Eac+VBJJGmr5OvzjA+6m4Ywj3p9zSbQ+hoR7hAkEXHcOjO7LnHFo1ELiPxiibJd++ZrmUQduGk9q
HnJpc+Ftk6Oe/v51GScTFjQtzwqXjOmDfBnrMaOWdQSIb4Gsq3jPzJlyvSiQisADoyn/uqOOejGN
6yT9YxOoWBPv+mf2Gjf0HjRwMXvhTeUXn6gQrm7X/DNDkJxnZ0ZirKOI8FOUUEUbUbW/InUAs2wx
AHlWgzUNE5b+qgL0yNH0VWGohgFmRAOjJsfe0od5fvLzQl1PzdDF/LmzY/FKJpFclteqSKynwTgs
lphpdOxmgsA86CXlzw8O/QxVTXRFylzjYQGsJRqNKeVLM11diSmUuCYjhvUFwTjDsPVaH2G6VDJa
tN0k75ZropET7ert3jeStfYpKvAgYZWuQMmJi/YXBKC3HnjQtpmLKmKP+tBR1fikruyzH4RgNnpO
lwB0IFMky21jwanWYKVBtKJOiVleSjq35ntRboDSmYuYSwsiOqFFsJrTr0vkT7VqQDekr7bp6XRc
uPHYB031VryE6h1uQonvLtmux9Lewjpge16YuYl7m1gEYdjwah4NkFi4ypRx1OypUBH4qgQvXUq9
6jMLDfba4xPlHhRWvjOY/OxvguOfGf+r9G78eFa9Y+Wie4kJDmUo/liyphijxSsgAGwYMVJJ+0We
d/ES9mvK9elCCPgyRbaGi05ikz6UVEBsjHSAoa1MaHpVXL8AMCjiLAdtP1Po5yiyyoQwoAEfkVfC
UtF7uOb3iBQPyt8A5Mp7tqMzwjgrOcHJc9zL3P4xFlyeD4X2OltRHo7eodBwAXQ5mpJEiitaNEe2
vPuLeA8+1S6qWH6xyEaVm5T1dTBkItBjyLLMGHeD79WebQX4F9YAIMYo9eOYW8xJnfJCw/mGk5mU
RbotEYmMcRwrDQerzd0Nvl1ZmpC1q6ZJ3ZKwe3yHJ2cugBEq/hd1JNJ7mF8So8ohMnprsdbWW3qM
Qu16ot3IUkYpy4N1MR7S6yOpqfJ3/moLO+hgywq9ZqRRzS3G4wsqqoQZM+FyKhj1izt87cKuUWt0
zl1Yo19TA5z8ZjU3pdzE1G2kEDerk2lEOtukIeP9G/KTZLMRqIomH3bhBq+s9b9RmBj5//r+BAZU
ongBkjz1AHRgANLJMx1JoQ2/g/jPLBOSfPdizcaaqySxRInts74ZU0/VLVK09MWRn0FM6bPYXxyY
fSazdJs48meoLDyuKfM9nXiaLAByipCuQ1ro3p6yAP65WqY+ThSwj3pW4L3/iFYO6HL5eF2z6pXl
xhm/vqiPdELvB4GlSjBfhVCDikNqauaWKh97TbX1R8ZU7VV+UNjkVfegPJNv7CVOmbqIdTGvhlgG
2Nq0OiLMyTPhPUZs4cIJXnn+OrE1gGzsVLLsoSSaGY0/P4H+RDGzx87y2e/8xLxTZDey03++E0Gl
Jk/ICKt0ZVaUzgVaLvtlepJw6MwUFwpk5Z7l3/93NZlCkSESxPjMn2gOEmYF+ciAeKiBYT58l0bV
aYeeGKhMF2t/5OmsZBELJZjKkqepbbioRczzHY3/GJv1qF6BEwDu7P+dmldYAZlpR4B3TNIawIa/
mKLP9fGoA656Q5PQAjtuiAK5Yx21mkH3wUgunRUN1CaMSopH8yg1z0CMkHPm8gLpVuwAlT1X9m6O
2JYlcJ5mWVGocX0ur/AYVwGIc43mVkZBu+FnaAqpIW5TkOYoSxYUJOyoxiSrp5Bwu5E43rxywYbM
qBViIAbolSsGvBWZ8YRSMXYLgLmM82KeUJYyjkYrM7Z6kzerkjTT0hU3PZGt8+S/rMLeyIY/HLkB
QWJIbA4ikl+6mXwHHSaXR7rZeFm8M27wl50vNtlHyW1sMaMOHnMulh+SoNsiIRw4xwpuENZhOOcN
IIi95Zdj8Y7WgydqWcbVaoAmxkhOE9/EzTyzPhCGDZC0pLyrBfsFDJyxomVTLRMuCVkLd3xVH2iA
3ODiAh0Mn4lSfuJ4HaJzPtVHykWmr/qP9YVxkugsxTOdWmHGb733zMspt0nqKLUeCOpY+mSOLs1R
IQeoPXwpXMvEIUR1Gol3oGozz4DhHPFZZuHdCmOoRj1Zq8Qd+p09e0vyGh+pB1fuM4SrSy2o99Of
//qE+kQHnzKLDkDtHJc8S6RwqguGW0IznW66jG6gl0AbulFcu1po5jUZ6Rvgh6iYHtLyw7AiGBoP
qPYmQpWm990ByqyM1PRXouKkxlOQm4MnFCEceFafLHK0Wuk4PTtsG8RLEI5PF+eZGKKyJOi0F3LW
rrVShQkQ990QABEJfROxbHrwB4UFNmyHVuG1NCnBIMswge18FnvDhS2UZErJY6kFMQH3yW4DEdZX
0K9jn3US2psEQI/t0+F972aHB94kYvwCI6rAcJJGQ17D7xmtBKrdK3fTjkG4WnqZHfhHpLH2x36S
S3qUgQH9ibpt5RqUDOLM7iXJvvpPLNoap+kSkD03QGWCCxUVbckMfdsol8TR2uXNwEA8R7u534Vp
/ouqMDhnURSkFzlHB/+PnNncwfSqC763YMq80+ugbctAsfE4MxPU9UftMmKAvMHEAJhqFtQ04Xh6
K5oA9+79oo2W09pBCCAt9KLWdytSPzjBOZgYXIFTG6DbqJy+vPtO6OEtEdkDuaTM4CfZCRzHyZnA
xzzp7x5WS3CQ/GnDAwODq/dRBUgOj9Ssft5AqYY5C4z3mdI3LCbNx8QrbCAgDW2nPgt/hwtmcNr7
upNFpCb7KsPCPcBia9fmys8HMJMArHCe4t6+5xiCtdR09l7TZFJ7HZaTEnl+/urtPvbHVEOxjGOK
z4UEiYxTlJFTVwUjwx+8Oh7/cq8lBsnla9lUlyJxt1nEMNn8QoFvC4PMl7SO+zvY/VXRj0Z7X2Xe
2KngD9OCPjb3gtDtesZl98bzzXmd5ysp28py6XQFyxdhAS/WWM5bA2rMgJz/mqRpbcviwvSayb+V
N6VcRGAFxWy8EjqTQPO6E32IfHJQCsLx0O+x/MRnJlyx1KpaU90ABdNJgHh0INgzPS5OBff0/Tqc
c8IrrKKTbWmtDs6oMW/ivoGPV4tecknV/o6J6zYc9vzuN/dfAFVD+8A1P4ZLGYMp7NQHgg0k37u5
dn6RDP38mVcnHJJWr+r3xjfP+joq5HDgkvRTz0qPBUCGvbZooxipbeUYr+ivC6PpIbsR/wfie89n
Ar0MKL1Fgg/IEL1gkbc81duTFNKDsEiS80G/NHIDDCUxpaczczKCKnwbgkNUDjSiUlMBdNXcaIe7
cceAFAhkgclKCLdKnefVsppL0zFxk/+teukId79j72KFCY8kVNpbnIhKATqHI68tRmjB0jpcxP1Y
MNqhiEPMdzVdZrrpzQ2YUmSfUnYq/bDsCWjYVD6NVzQWZWzF2vaAXSXe0fSGZa++vjqfCeyRZLV2
JSoGyAnqamMBs/KTlj2B7BS5CpTTjZ6hf2iXvXBoxZm3DBMEEhHfiZPNE10eQzZ0kbvqmKENXUPn
eZdRvBEHnPEmK+Nv2PBePKlJgZl1wUTfro3zrW3kgx6swbXdyfEQzUHi4BMU19LGqJkJdPbVVqDf
nC16ny4Ba+r1RL5/X6S7z5t5fUNj90wGqK2Engd4jZ94bz1SNG9hELpQjcfCK0PIUtd9XkMZP7UM
ddtlPT3NimdTQAD0VrHbBZtE4EnP3Bae/WVDkEWuelVXZ+eCY4BlVFc/s/1X6GG00MRG4I9l1+Y4
G3FFJJIfDyZ+Iyp9b0++pCbnikOiVZRExCAsvny9eBTNe7hlXmDfFw7+Ccbpw6ld3P2+IL7Lplcz
1F6RGW8eWWod/bTLcsdLivRdl8Rd0XWIsv6cl8wOxZjms3ltQlNgWAg65a8SAeWRi3z01CFEnM8V
ti2PnYjWezOvqGJFmD0nm09jImJk0Z9Idp2dsjqgkVuPfVX+IuteXZd0gewa/C4jCpU2DSCdOOrz
5N6SXPX4/6HHScOwU5/pM7F/oRM9DwGxQstvRVenB3ym49mC/jYC0SkQgd/onBFfc6+6Pe5gimo+
YQGdaBddAxN9F0RiMMBbXz4oB414xBPFiZk9jXmiV3u1Ob+lEZfGK7Z8KuTNa+UM5iHAHS1Tj6OJ
ZI79hyRWjIUYwf+FNL4pt253VLgZtEoLWGuDKNsdFZ8cWlhEDx5LtvFLB6p00HS3yqK+MuHUeWgt
rm8Xzy4rrfX31IgPsQCIJ0BsRVxgjRFub65R1H4oYFFDCv7dXSmt7toRvZaN9rsWtGNF17eI/qPC
o4E+Q6K29zRhUKIDL+Cgw0cip++Lbcn5ulxSVJnZzsyiW2aUANH7MHJRsh0hXHq9xiJQEsiRNVka
XqsFU0c4DyTeZfFM8RcewM6igXo+7Oecgb5rdWoHZbeHAJ8g4WICN6imQuAJCrtP1IqY5qenxyg0
7ByoIwtvt6k9cA2ebFukqNrY46PpzzZ3p1CCHDj3pM265HnvqbX3extaLDLcEf2xUFSFs5ZQk2Yx
w/JGlcym1/5JRyCRSan5hZJeePODhSybt/6mgeLyPQsheEujPjqUhigPBcvoH/Znrr6XKdwei5em
lgA3Atz30aufw52tgu/Ehwq3lu6SZAFTEn3H20d4nJGmyymItKsB0xk+T/whiiVb/lszzt6toWc+
npVqFeTN6PRTWHkp4nAzpNC7J3BeixcLSPQBrH1rpYbsylxRTTXmbO0A8QCuppaKJsHYckLMR7QE
CcrYnn9UYzVfIp133s6wLElad9bWXGw8hf3I3lNOdw4bPIBCRkAHYA4odyGXaSRryQ4ngD0iiqaN
v4uOv3VPvnQUghqCcqx2ZBDRrKGII9YV8G1mJxL+jUNk+pOnsmoXCKmD0/ELCNO45/n2kKhAkqS1
dXyjWwenZxitsUdiGfPWlnkzewWdDLBjpEWOobl9vwL8HHMlW0JQP2zWIcNCuHkUYwp7Z2TVRhWc
0nB4jktt7J+Dp1FK//ouf3TYbGvPEoKHLsJTXAzhCpn34HZN2pJtV3c+/rMHUVMKqMaa4rleaIdy
t8/lWEjK+56DOUE7VFOtBmtGans4QUHjnVaOZ9+CH0lFUn+YcgnONBEUxWKxzVDg4JvjCTWNlIpf
vB1GRZ6N3dJWoU12K2DAj1E+Dr+E5vBIowGYY2eTChSU+nGTgKxXB2gHKFeA3xZ53qnZbbdfcJj3
k3E3hWluCUznAy0/JybIySEfOK5JljuaXpbyDPl8E6645BX8RDcskMWDtFqmoE7ATfHTkYCRBQgX
vxpJyv5+jWEEXRq7qQj4J9ggD0b+JCgUo4wtV5fKaagMHOcr3VN62cU+r5vg8T3ySDugo+MHMkEx
GiznhkZAoFpcADqgKJtAVTmU2v/NSNx2iQctCMzBY7asSZeXhy4f698AZP5LHntgCIt+kzStWtG6
z/9AG1eubAsFgSOhUqPIWM2ip2gV92jnMoLQQKPbOWT0melI0mBd3epYifDX5tzvIw+/bgrog8Xm
eOQqWYiq8KXZnGKpUSCOXGLlD/b0UqtZ5DPhFTWoVZvwwCWudHSXNFylJybJpms+JK8d8VDhxCVe
QQTxvYoHhoOOdk7ngcm+NhkQlltXJBuK65KVEfD/l+wW4atAUQvct6DplKl+PgpkEwq4ac2hHcp6
rQJ2NucAtuUhkmcZKE5IaLmsLqRsoi38+z3LSqQdknVEGXBnjk3BldI60J3eYANWQe6pZQooazfc
Cqht+Pny2q9vCPhvidAdfhTed5agqjIbfnzlfHIpiPf5o0715UVQ/ncSEPU0VB5as919533oS4lt
/UaGRFIiE2EJLbsh4yW5rwvqV1nl1Hhex9u8E8++68cGw6Kn/1PzSaUSOfOA8k/10UpyL+UhycZ4
QG89aH3wYB42kYaTe5Pt3Uca6SuL1xQ+VwkYPrxbrQhjfEKB39cUmI3IWIKIIOVIsoFk2KpWjA0S
xOzmR/V6LaJW2I8sAPIZdnTlX0yhaUN3zOHYVTyxSZIez6/8C7oNaLSsJOXu+mwgiyk9Xf9vrZ+8
JCyHsTjHInCkBO+WLlDBEwDi1gNyPoaZpF4VXJ5JTtpLrJ6CJCRgfoJq+kOjK0IgZK1B0+hoo/s8
q199tPrQ75tCqBe9d5Ss9CCGtxitG+ZwvPN1T3BsVPHhyzgR0pPp++qgIMNafGLqY89QzQYtZC0y
kRhaudrEFRwJaqsvYlPbtylao6q4AdLH75OwmRXAsIqlGxQ500duaSzSdIaEK72p0jOe+j1i9ysE
fptX4jVoo9kaGzehhOP8+xA8yN7SfgmfrHpr8acS+u6sCVmvhgn+n2rHcJq3KJxMPAkxp7yY1Xbm
/yRLdONtn4fndm4upWNdDUWHwJr2UdM1tBQ97d3dCiJobMkX293haGovVz2R1BDrK72BVKpA4STf
ner1Ec5EBxH7yDIDtcDhqmsLIRcJ85EUtAD6wNO1xB4QPDscyvrXxgjYzHw+hxYEyRVdQzlNJU+W
UiokbKqE9B9ZPVUQzgcPZXCl3qSqYj9fwiakqgPtpof0Tx8Qa+BgI6dOo+cnsSIHP58dAEhqKfdb
jneHlDdtu7PAoA2xYFcBAjUginP2Gc+4nrZH+vrTxwpx8P8Ppp/izL5tNs3H+DhTOJxFQvoXkBSD
LsZD4njmnOEqYs5l0m+fu8nNX4kmTz0sPtm3SF3piYgDv1/kLVEd/6gjoY4BEg4UQTFRfSMf5Ubc
b/5i8NlJsxgH3wImO5+QLHhdG8wR8dbr5lnGGNNkoK/ooGOVJOe9cOm04SWKDWrtI0ZU33O+gXXk
Yl+QW5Q4PN+WQh02RYG1ZCq/Cp0t+BPGu+wcnsFZ6Owp3xpx95lQVlzT7+202oLQ40syHiDA+E0D
SJzT9P4/SZ4WXkUpma0ExaQr30FQe6UtJAyUsNqJH1oJnIYxWg6y6z7E0RN2SiIon2WqbySApBLW
HXTkcbOPSG9/u4sfM1kuRq3hXKzuaoBfGvSv88BtiPXh/FR50o+c1NFNarIpMJW8IW+iu5q67kAj
ACexjkFg3kJ++U0KIv13TDaXrY8udXT81mi1xUO3hFs+MrFIXQuUXirD5q5qJuOSlMFrLtlUkIzn
TyBCyShcSF+wZ8d6xTFnIXjgOQmaovMwuY/RIk6MaSr7KF7khDsRQ3Sde2Sgt/6u5sxhuxTqxfC2
JnQslb4FGd8weutp7xltGtIZhiWGsWzaLS0TCS3IMQEHflwHosQJKrqeBZYebtKKx/2/oYPme5Y7
oBcpDOEhDU/biC/Z4E+Qegp8Uc8bfAfLnadHtUJTJFBa7AdzeAttvLNwoR/aWFPEgLbMXM/Uh1Xx
UCO9xuPbeuC+uB0lyQKxSFg+tCaSgJQQFHvGWxRBN2uiVp4PLW7h4hGbz3HkbBp5sL/JrarA91yE
uFMyrDoLbriG3oArFT9xb2iXNXEcfufnF6OXP8YcuqYWUWVaO/wA1xnzx1uMIezbTFbAi86d0Bhs
C9nK4vK76/zPwl81hS7T6tWorNs9e/tb/TsY4qeD8sMNh+/0Q0X2zRdGNX8xU0wbzooB50KLqxiL
scmA004yDe2H+BTqn0tUUoVQvSrYw79gOc27t5LZm1CTloF4hPOAOVYH/VheNWIXuoP+QqhsanN2
gFUOz+HEwJa64FUhIsSjZ87Xv+8bv8WmRy29euJFNqAsYLBlVTkMykJb4f0OYr1qo9qBeX6Y82fR
MaIemCG3G4c5F+QG6FDkQdHj+JbiS9Rsqw8fVWwlzR5u5CNAGbqW//njJNDKAmv3V+fj3TUE1V76
7L8HJaJFR6TiXNIhQbt9lEQA3Dv7Yd6J0nJS9JOXTQwyiF1lh/TJgUGbPS1w3zq61Sd7doFa79g5
2QwOdq2z8Rdhgqh9561z7YKT6nyNQ32Kk0KQsnZhZop5ScfKDcwskR21gDwq+/SYp5C1x6PCmJc1
a98oFQp34koXPQtjmETJRxBi4JyNssIa/4mBkzIShlNcU9y1j2MHSlobxQYiTs5nGx/KWBdeX/hn
KlcXmhAjctsHjD9k66Jt9kzgzm4nSpI/IGLDRLFsk/1UFIO1GvaR8vKNeRNRuEN+CpIqLAG0NuLU
Ozbnsx5Md+gex/bueMzJCrUZz1swS7dB0rAdp+eZMcscnKXfaxpa9y/293f4EEgrOw4mjFNZJ3G0
RnWiFxnmX4a33S67haoe8OFEAWtpq5iN83gEUelUzZmPHHfo7/LCnuI5ozbCdnVCI3gdzgGvyIJ7
ohjkFeyjS1wvYq6rpwReYsajfv9PTQo6TNzn1rhD9OFnZRXD7U6zbeCufg6YEeGR23SGuxx+rrgU
G1Xo7D2P+iKVA5cN+xt2QDfgruzWpthFgcBQqUMmj4x0OfkA1AK0k/u2co7UZi6KxOpxYreGNHxR
4EiIsnLFXGGYaiiogRDU4T/bcbsmopXKPEvj5JkEj5Uowu4YJClMgLqh/pyHUeW7x46+LPMdrA19
aNpVgTa+3y4eUIIDtO6VC8f3FyPTqoJNWi9IkA6UbVt+WiQ91HpHdOOuXlE9SSEETRYLONPzrx5H
QpjHsUPgQE6tpfMmjZ1hQl+hjXNI4J5pCddNRpChc43qALaCZvxBqX/kGzeTa2c/SKpRW8Rxrqax
Gx6rEWd8QxZJuOA3bHaROmEmNi2J2KZQM9QLc+grWH80HhjGXgke0xsK+NfemUXd/7Ocs6E1BO0y
nHdNrFczxzG73HtldjDFTI+H/eAcBrCrSTIc2xjcIWKAhvbNVF/6gGLygv1kgR4zEtpDq6ami5D2
9UFtO2IeyZuO2IOaR36cXKYyhp8HcAdxTe03inuUPjZtWSj2Ab0cxtMtnAjpOHfR943sgTrVcen3
MEHYvyRLvymOiwvgmUSjvfM1xK/g3Mu9PXLzehHUNpyUr5foqAhDg/rqEMJHHnECyF8N7f6ic2vr
EFQ3lyEGme7aTSdFZ3udkAgDeSDtv9ascP4Ug4hJj07o/4X3mg0QuPA71pOA5Q+G94uDlwL9533a
Nfy+WK5cEL50cL3wTt9oqw7HtDcgKu6foPl6T95rZSaesFBQ40Fm7yhVqo8V8rFMvBdNojgEY1yd
Bf288um0v01lhmHEJjvwveIhu9+xMvpdhFDSrm0rVqRMP/ZrrY8g8sey8Z5aReu9RZ2ZyxUicfYp
mkU2aFvxjOmXn+wn2X79ZCG/wP9quHOB/ky0cT5nVN45US4F11HFgOdLRP4n+HCrwlMxSelbsqvi
9ISLvFJB7LQ7fW+Bz6wLsglmZ+YYNJYWeHLr1+RoUhla5Et+fjUHk3/WHtgUR/8TMywQ3DqGIInx
UIDUx2Ybi8jSnR8jd9RbX7JSV6VgunesOc56jR60vPTuPpHOATi0JNmHjmI/2eYyM0/v6EcAZDht
w1G/oqgAGAANOqc8IjHZH7yzbY43HmSMbcnGTs5iODaGCMMn+XKv/RZIx9H89y436iB4f81XoQ1F
cKOoLt9H08skJOOBNDIJKUteFI7xqHWZrcFfq2BJHzNqeAw4g8uls55sz/udXHmYfl2F42EjA4al
JQ5o/UVu1Iyb7d7YqE4YNTcE1M2iQp5p45+gy4smwrLUBM6ln9YawNROQLQKpA8v39onNIqUqqS4
2QOJfR6obk4QQYJ+2Zy4TVwh49EZVM2dNgdZeTPMKirMz03tY9mWVJJQ/U28dulciAU9Rto+CFYv
S6tDedNvg+04AmX13IymUFb1XDtYV0xMKnTXO1N1oediIlyyWwQBf5QVOW74NuwXVnxq18bdhXrN
SarBE7003lGKRtyraiYn27eRcziK4QH97ZFrpvfNqR78C+B8xyNQd5+DkjOBZiVpWpgaJYAw+hpi
6Le5sNpU7HFrBEjM7jKJ+jqoxvhW7IFCyOHJB6U/gqO/gk1qiinf50h/fu61d61ZjRG6dIQsK1ip
xr1hDj8Dyn6YiAWXrUu865BtthljtLMdG9fHabSsSeMSDaQhnoiyG5uVxyyyCp7z8g7yZt1w74BF
c6ggGtlnXf7bZG35+g60iVvTDtao9EzBKzM5z8CHVSEVqb2M3SlzsljQnIJQbPaoZpXZUtWAcft+
u0if8HI9zfR3VzYfevKHXNCBnyAL2Q==
`protect end_protected
