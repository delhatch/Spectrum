-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kFVucXVUnYSKhVjoMsK4xdHFaaEx/NijjeNxFosi/yiTomqF8LI8DPWHkAuMOOhVXu64Y6+0j2lo
wX8sxOVNecJpge0chTNLa773ajsvJ+lvxHBd3Hgxuc0GNiayTsE4D49ZM9SYoKVWETvgU7r+COXe
ZEUlQyOcCcwQbR8Cidi2YYgqbj1BH60xIxqXl/TplQabKTQy+K3j8TJ/RvQoamz2bxsKIvDC8YII
KUkATS1enm/+xpQ4NSRIiQZHOm9I2DEyWLwhHxXnpdNaPnpjdhM81m0nm69kyoiiLQAuTB0d63QK
NF3yt1Zaj26l5vfu2Qwhlxz1jMTWyxn7cxxwDQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
ejQYKDb7SYS0at/9H00pTmzOeuBIzaK0iuUxi0iTIiAiUN6IxB2g5HrVD9SH7cIne6DgDqdMP0Ed
UwYzLvoLu+HABfV7ZgEXNzQL9M5di79DoIrA9wtr71qAfV/FzKD39m03TVQvMa0fdCTmjAg8XMrX
NatG9NwrmmG6jmayBJndzyzrx0Mv6M80GEaTppAPg4Z3o3Yf8HkWsBvc3DxBiBloLzAaaHP9LkIu
Q+u/0mYXdLseifq50w9KTB/XA7MWhmPrWTVIrIqS9HcFEfPMhBDLl0U6oFtoXT4Perw5XWNwC/VQ
eWJiNm9JLMsS1b2bUX5CoUVPy95O+v5aDFxayRBMwng6jiQlEUFq2mCITlKF9g0DPGR6rVEI43eF
30pHUuJqTJ0Fa/EPZUrj5x+9x3bJoc1M6xl1Vk+40gpSZqTnOVpX2QZQemZXoTu9QdsjJyhHMN2Q
7HdqW3MjM3QT18tqviI2zn57lFTWUPHv79jHSKLQF5x6ZDJEtl0fm40peHFh1YVm8wrtwW8gDMNg
i7xzB0Xx2xhOg2wXXgKYQQlzmK6umoMkmtSnmgE+RGvcEZOlp+L8U10muzPoa6zfw887HH/xsCGS
OEKR9etbZ3v7lGn/55WjNpWgCocYE+jFGwhw/bdiVh3XeIJrhiRRvxLnJ33ZneBdUbKXXri5+pvz
UTZCjGfb4oHnxKP98f/2Jkqm/Gv7sUmjsBWIqLGi4n0HXQ84UJrLMaa9otfFRkVhrd9YhQJ3M1/m
GLYIyFm9Q7RW5++ixlcZwkUjNDmlQA/FPHFujae0lK+xR9JSxZmuCEKCYqWjs/iSyFpprA4cMSbu
Dnqd/8xYHJ2o6uBNfdRBmEhj89s8WN3wVk/LlAa+fJvb3YQ/vA1fbRrXNYwajPw45MT83OE3YrNn
JrvuC3NfiXswrOot+zyRetDNHPV6fwlTaYOIIQdQIXz5ZGbKRteCoUMPwkMsqipBAsybMqIIvaO8
FiZWaBRH/7n7oAtvGYiNKaixmMRaCfNxnYEwCPkPajZ/8ENhbSPLJhB4Jf7qwduPvT7wXxsgXQRb
sXB8F/LGe1m+9PUyQvlg3H2TU3p5JAAIHPfM5YYSI7U0EVwFBHVbjhVaimlAiLZiEwV2TDtxRw3M
Q03iZXhi/kBFKdgtWYDHbP4o9UXCiydmc7ygfojQrVwIuJq/VCSP2XZ218UbGUyq56O4E2Bvo2Yt
GnTccIdcF1E5a/aoSBpHUb6qkcnX9O4U3Xu6pBP9xV6FK3uI4fRA8U3P5CPLuqwUoO9292cW7HIM
lmnuY13ztidwxBVXqqNVIrWe7mS1VYoYc5DXLiVCb4avgMAWi9Ri1voa+0YXRE2IPngX/bk0HQjW
3rtBpoQAQya2W92XymlJynb7DfvKT37wIF1naHVMZJDYsAB4EFlrcRdOlipuH9B2iX7XZ7Gi4tMp
zohWOwllayjCEWqsJBLweVDlYNMM5DxAluU2v83OgPt9Pt0NK7OKnhwdk2qYX11fJEmGzmep5Wkg
DAE1GqubyHKb0ghQpNZx0qa4QLLroKSpC5DApr5lNdEM0fyMps+y7EaqRbiZ3zxaCHzjv/5Q5cQ/
cHrt9snlXLHtLigl9u61Kp9Wne+K0a8PtOdTehIINybl55QqJLo3cF1V3MmhMU52JmIOIg+DhnsD
i2tn3y+vfqYXg+FNiLFAt9etAQ3EKQxaoBN60mRkwtYHIkh6Jvj+4dSSKOS8N3N1IgenGSgmRbPJ
hIjbCpicXST98Caqbk9w3YtwtV8XgTYgYqrn8+GRKrjHU4krETI5YJspMYTnsXUhEdtWg1HeEzyz
tX/dEu5g5wBZntr+WtgbBBD4MIrJqdsMzHzfkCmewsOih/wb6M0FrFZhKe40Rxsp4nziakvlFahl
zXDuntCa2tmqsYojtA9ycvJGxzrMF3+3U3RHaVeVyNHs4M7OPMaahQtTHQnR33BXjXHXtHXsANkM
d4WqzmD5MmqhRTQ4RU7tfDluJpBvDW9A4/RXPFpFl2bvppLatBGMXOU0jK/v0SOiRXhnmI2yyF46
H3KW1kEiNdm/yp8t/Bpa4QWtFu/+90slOgWOzuHALxCE+tTBcMC3j5qNY2SoVwsx/ufyMY5hjke5
VHCXcPCKdfMnoU9IYXW7GI0p0x+Y6AS8NjwBHqURlJ7EWuGXGmGG+4OQB/zcvEr2pzo8ImVTUBfA
4htXRvJhkSWTuxNOZKjbbd3rwUyeFdJorDv+OLqtclqsmwWao3xx9XYWeVpGrivYBbD20465B4IF
YXCyuAPnY7GhuFRgb+ICDBgo9es+negSqNPCe2a4PDYGiiZbvujxzWIlYwve/GCZ1wE3Dzn8Au4/
4gaKDiXp3YmIs5lI4j2KRt28ACKlNcHZpOuMBfqDR4PNwWC2zCFCgmYs56H1kYa37MFnLxvWdqFG
k1cjmf//qVvIuR56nQXOzxoj1Jgp/JBsLgaAgBdXhzcVqZUNgMFMfFEuassxiADWNQQMufop8CVP
+zlTNh0VmoHjsaCqEpp4TU6CG5Xn2Hx5nsiIoeWoChNjFf8b6E5cuJviaHpJ9WVMq9lZ7mrHWINs
SUp8APODaiwoQp/WEYD2hE70+BclC1dVTu1OkDOuOTSr6+t0Y9GODK6Z809dN+iK2ePJ2/YPehjq
0n9J/2S9cYVzdZt+tuCKCvfTK6xT6/km3U2joBRCnxmlo0bWM4HRdKg0yS+uFzL8h+empXUX4+Ff
AeT5CxbsNrad9hsNchIcjK9uHuhd1VDL93gceJhMjyqe1ZMEHJ38cweC5bIVfqfcNvmT47IHXo0v
M4IC3RpNmt+DRonwGSi2PldOUAE+rEo3Ovyc840TwP4X1JaSDjnn+mX+KCV4HTIbxsZGfeK94sjd
7iRIvMTu4banF1mqVSJYra3ptTS1P0U1/9AAAlvPWfODRG7ey/x0k3Hf/7ucCYiKmLWMaqvxyuwB
YoD9MtK88N34htkyuNh3u1pJC7r0+CX8Gf8FKWYO1zpMHVx+gjXr7m/Plyq4F+Z25qz+MDq/uFHL
7HIEIbg+x1RHNczrci5HbiXJHVlvEaTCP3abfjK2VEYgAHEjQoqgsLJat4qvJtm2PALVYAbJO4Ix
0Gx0GIWPYxHh5PJNA7kJ3Y5XXVodeFXZqywAHQQyLCfBek+UDRmeDqrGReCarSzGnjXdiHdN2RpD
hmYk/eHC/L0yideyImAVTG4ubFrSM/MkzfN1YWGmOjG3NFJQstmqpipJHojyyUlQ333vg8cpaiJL
BR0WlLu/B3g+uOlpyUgJIbTen4Q0TBCeW+BNHg7zRQUD9YlsGeTRRqqzMeobhr8q/GmfR8LlcadT
TNMfmYGan5xkY0k7AmCx+U9qW9WQ7MkcfObPm31mkataMOPeGRGR21fb8hcX6Z+pDPTWvBMkIw7A
t76qUouJuEC1a2Q/hHd4Lx5HBjEKD9KILmp2BnKNYa44278rtMasTNqshDZafNrCnjB71FMJD7Ob
v3JgvYDGczZ77DXLik0rFXHnywqkXztRFQt0QB+iq31gPWXsIYkDWGFYqU5+aQNJrjk/CP0i2vku
PytoMF/DsRYJqwfXIpswJkuKHsywQRfPLEh3O0AApaHuOO8vmggC0WY+cLGm31MUBA6wLAe5o4BZ
zm3l8YV+9Y/uo37tgsK1bcc8p6Lta0qauYDAtXaPVxJ8Gzcpa3Tpcl/EEJ804IO9wDrriUVIQdqC
/41b1DOH6VoFHdyHiErARmL+aue97NLrTW7UwuBQGfJ2lEJhzCgqCtX/MmCfWthN3jCNdSD9ou4M
jyPlqa7gRHqZk8XEx9TAEq8AlZCcCA//Ag/5ULN/vm7v7DmeGa8l5dSsCfccrcXe5mw8kajW0VbK
/Zc4Dun7Av04fa/5Q+PKFDW0ySw9l7XGpsI8Ej85i//wnHKmu9EPb2O8FOzEXRQ3pBaGm3oPC5O4
8EA+5079u16ODvHLEU0ZCfz1VYiMaUfbf8+JgUGSmDWkqq02oCLnh5amKpnXeh6OVgS1GRmtoRXa
rqTWdZMkYmVQDpCVTS08PrpKS+Pny9K/u2U6P9R+++XAigruk2WsXXt7YQ/Sl+SNTzVLV4kv1185
DKGhYXORsNH/uQBBW0VO73xYZSqYFTInofbMQ4PTKag3n1UXLWyYxg0nKscWbgwAfjUOioMmpT3m
x9boa428eef6B/dZBKe/+HhPc2EhqwuRDi0gNAx8662Rmv7wedsZLdRhVV/w/TlVv69h7Bz3i1TT
O8ZrU6hWamhOToQJdheQjkzu5h8xMkSIXm6z1YljIoaELsup9V3peG8MwTh4y/l76S4KNhvxk4Lm
M3FKNQyMW72wKIogzIkq7p6YfbmAk4WUJbNgPFXrDIEp+RGBx/f8KsMjdOEme1Fwg3c1MB2KCI5x
6iCQeIaiSlIF2qDN1UikW0EGO2s2uSoVgPxsFhJTvKZKYcFpIDPBOEkJ96m9CrFuNwew0gDS7UVK
IxeyiKZhY46sXjTlUHNc4HVjp45HJJTw+t6nDQwz2P1eqBXijyXc/1/DHOSw6UuAIzXVEsXK6H94
3R+ZsDfEx1rBlKANkEnS584k1Mmkn9Sz+GNkTWD1vrhdH129FEfJvLYdWwVcW3X8E0apYxAjLui3
kDbg7u1WYe3QdW31pZ8KdNR8ZLUE6ReC99QqFN3dIZrvRJ9rIYFLPOl1LYW6Q3l7x+KR0oWayksx
GT2fTXy3Smsnh/tfVOe55PFMuZ0jXPqD3YG/tI29Wnf4g7vZI3ZgM+RfEBGoV0wmN3KSlTRPDX+W
Dss4I1DkPzjYUbajp0CbXRVCGiTnGKpV09RUsf+TOKssTzO4WGGmKEOepKVp3230cHkfVU39HuPa
z/50istKfZVhjq3lvSvkJoPQjfibxCQbFNcUyLJXp8fpbAlgmqCtaXZKhgdtPJu0hmgb8o2cu1ba
3qkqRf9JZ9FIfQ57t8MZWjDFm5b366jwk6JmA3lkOO3TeikrqBGsLO0V4k1U247pAiFuJAAv/JRv
R6sAiWbJImZopk+QExuEdI3HSOJnoUKRSnQgpc9cNXlpa7UAzA6jMWYQfbYV1X7m73AcKVprdFAh
ivAZ1IIgMMVihTXN7pqU0Ew9mEAkSzQDDMPW71488RcsoUVnN77+iFdBBKox5R2/zm43iEbRkyf4
tIVF/eKjqacGtVNttcfKZGesHykOgUpiyC0GE9ABylMroxg2x5nkn9v6OVxuWDVpovE+weLyt8ek
A3FuzeAvZBmD81VHU1kjV6JEeOMbql3QZjRO0hh23tvpnrJA/4cEuDGqZyL4dFvh231xLQ/E7sHy
ZTUvdlUBfNqLL54YyzzItR5lVJm16nDkLkiwHfblChkzVjTNrwmuN2Evii/UOLugj7kST1nmDCac
usCL2QOXz0banbL9zqxL3GFLZjvj2Hiz5k/l1zeYhSXuP4+eS35v0s9JKEO7o+dKasUFQ4K1noEr
bJCAcMPMaU7iv1N5qiWx4VWVjTAXbWlFucXLZfIj3YCnliXO8E0ugMpKdb3NpJxSqdXB51VTijzq
TUNlIu80j1semT/l/Gq7g9XsjyErLTq5Vx9Q5rdcsgcdMFXBX4WMm6XnHaz+lRp2LIhpSHlUIlhw
lAWKC7AKqQoqbEapufbPvu8FPonpmgtXyxSnD6moFgFqmwY1HigV1YTkuH3wPDbbUXCzl4LEw9LS
x6BE56qgRLPZzKBcCGZgtJ4t6FyXGH9rvhUjl8B7L4CvBJR4gjVIFuRfy2InrTaGti7ZBV1UKiNF
SQiXpkuDXdyzyUqvMaGDiWXONnJfEe3myxVS6bICh2wXICcfll4XnhMFFD+TMkbjkE9Y1pbQTkVn
y3oCZbRqEnTTULGh0TRq2VbW/IcYL14cBLVZbQKmF75t5ThYr9GXWILeUU/V7XzNeayh/6LWWNMc
hKvHbbFQlBCsvwn1rkWV3ADT8FFOjZTeygGA4B1eDgQFnGPnA+aTSRUxlLcesY9g+KY78JoDwj92
041jE/G7KlmSQ4SWhT9lsZjzcxrBBiuZ4eNnNBMRl0x8oR1FKqLf+LYzRDkWLR377EM1aqOxkJD0
LQ/q1Z+eELFDAUudJNRK75T0HJdmv1HHYrN+JbsddlSIUlOZshhRy6cpunQeddJ4vqCrXBMA9aYS
B/8YvvVe4lc0GLX9Yct4a173Fp0KtOJxul7WGX6E/nKlmr+cPzu2Gc8QzJz6o63fA1GiwATP4tcf
rCvVklju+Vm3MNffJR1zFpLVnE1yXL9GDkExxJXRlco+jQ7xObPBUSwuTMzpetu5oas9W/WIAlFh
VgE9XhM769RHjvjipXGTQTBF4t/BAgR7GfOkNjxi6tADI299GjKfy95Ih68kRF5X4rVpSM/EU0M4
JQMKfKJkrf2xU6DizdL1OWey2glMj+Q4Cw28RzXLL2YFhiMcF6yopChry0pqjNdIlxO+mUxlc0e6
kz4goFglAiBpAdLE0gWCt9oJlFKkw6Ehq9PTyidiYAiMNUBezWAXSqCYyVZ0Ne+xRJrkjY84efp4
EromLgCAfdfFy4G/x0KhcRFC5zw0Im5tmbTjLURdy+qlsYR/OyUkvWcVsX7vScWj9b+/bYZN2Wui
58aneS1ruN+PcQb8tVMfpyaQuGkS2FlPHIRu7fhLfJw/urTWCE2ByJnRela44wEzyx4eSZnA0BhR
4GmX426dJf9yz4Yk2ak/gm9rdvLcm2vVKRrTU/XGKMds+qtR6/SyrtnyIS1FJ8FLkONbmuzkzq+X
3tUYJFRWEnGwL2QVOeTpDQc68cCW8piCGUO9u/gURMrbCooiZ2DAaAVYV6x3XeJa/lKPWBizeXah
b2wuGOwSdOD99rgK+XPUY2EVVPR/cprb5fnDO026lSZko8Osq44eZuuNr8uzLx5q3CIPq3QQhrnt
0XjufdM0tjDAqT0WKq380ZPj8EydrAxFgnjizUt2q8zp3v5a0dDhc2urhXXusYxFqZ7LKKDiGVXs
YPM20Dt4jlww7M+Xs8YUnhgFPAIHvHiDIVDHqXgq0wl5VisgQ907+bvKU/AwpvvrxoJC5RGQAC9+
MLXWXaO+DtIMbgZI2TewmGtZZl+p/WPo1fXKDx4oZb2LklSNcFUH3rYPzq/MMBRkacZPgsXMC9ZV
9IJY0Ml5lXrDiZmgAJD1gUWqClqWiyWvIMC86IN7Ty1T6Rch7P2Y8zmWx1sICWJcg+mvIBxYNUCD
QOVvGw5NAQdlSTKJ+BIjfzThMn9+X1b3r/2RvEHIDyU4msBxCyhnuguj+FRzjQjLLd99QZqDkput
ULAtj4CMj+x+AqQVBwrPGkQ7MvpwnTqYy8rfAKEsiCIe5cmKDpubMbBjJkiIkSNeUvVTrDSUqjlr
KDlCH1cNYcCh6PoSlJwjtgRY92KdkfGBXnuUIwlRqL+G4OePvq1JOh+nxsyPswE+STDSUl7cXm9u
ywc5MuAbvlj4SkKr+RVoq2Y/pKOAk6y/HdEQJuFM54XZggEuN23e/Jf0UugGvc0JmUlxoOuOcAon
N7I5sqN50WbzkapDoXXH2Ln+3SnOQoAfq1OH3MJ/gxHqn7UvpdeWbFtWnbhkAQlZ3DiZNcE3gLeq
ibsn9C3wpoKwnS2AFmzy/ig1L92563lRsRa15GEEppVHwuzdEtyBjdxbgjAJ/YkyYiBPYu2+uvh3
XvpNV7DeEx9Ten3+UHJUF+IShYj8vlsFT1u4sBuKk6espEeZnav6cGTJT59TBSPeIakpzvdTrJ1p
s9JYQmLm8MZiDSBEF4+73eXoA3+S1M6L1t+4MYWblEE9GYE9mXxKIMbzpBw/OClMD0uDlG6/4Sm6
QTlQNi5OA5eCRlBZdiNsSHykPX5x3zlsdaiI7mmhLVlIQcqHz9gavqQ6F+YSyQbcacxW2mP2d03D
18waN3fxvqekiPSAAIXYwifGB0Ok1pprYesDtWKkjR50Gn/ayUo+kaIP2u1IcMrU8mmmIlOhmN4/
ItwBMzvdjde1TiQhMZR3BmFhINCCnnfRcpRir4uOvBm4fR/EZo0kua+AyxpbCEztcnBJdDV3dpkc
OPFQGViiBFBJDAuEzyxXm/aImYjYFACCg32j7voA0T8t1rUdnXRnwbMWIXZyaErLjyrDnqO30ePG
yj0k4znN4NCsEhP7XEJbpUpq4cZQdemI4Ctt5cGZoeOh8EwPDfppkruqN6r5L77JJe1Pp1r/PuS8
pTE5L2DUJ9zK3NjHmjleCxYWtVeflOSu11LVUkm1yZQfvolpd95KAS1bgQ0YyQARCAAr+YOAZ60d
R+V8gZqObmyR2D36ONmzSSM2kpI3XI9UarQqcNxRArCi3YVyoPPOtQEAtzWZALR+VmO+px/jfBN/
pW/UuNY6sgVWueoaCQ1nOfBpyDKaI9YMxJ7rYUWYcyxHwqVYDG22TlP6lgLhBcCjMa7CjpQpP2ca
P19K0S4Qve1CYS1C3/yIGj0Ne16XLjgWWg2IcqqY/bVwQV9fLYll1M2D9vVusShR0Wr3jDqwQ4ft
exX0pYcyjWFwVxcUTQG8F68c3PPH02rSNMs65YDvLJRKLm7BOPEk+12mp3EmgqgfvstURWi3KHMo
XSv7FXK+X1m/N2nO9rL6BnXsXG/PnbdY7JlJaNSCDvD5KU1PAKcZ9IQ6EVW3sHLT95NNOSyjVz2S
Xjktb6BgEk0aJTexMEoaCVozzOt3NqoMcfVeb7lWH/AtdvqZJ/znK4fD8a7U4iOBHWEleGmkZw4k
bJiqDp+sxy1VjTh6jV8AzPLY15VHmgDLPfGE5CAX41r0lwhNhsDhrUCLfsVliFNq3Ijaf+zDfASz
OMptAzKT4NY9EX5srHdlwQ/ZiFKO28/pebR3iyUf7Gf/cqlSQ3ctpcNG3gu5aW8qczWdxtmxK9Zg
zOwaVgG3PXgcO747+4OmjP42/OnBccj0Zwwq9vES4j7IPFLgnXG/WTbWSuE0VrONvb0NbV4GKi8f
41oMD/nmI2UT1Ytny5uIXLfdzCoQ3hS+lN86/g75R/yGBiG7TIE7jaSeyWrthXtpUFhNGb5LCj4y
5Z2Zgc7MLuyweJNajF1NvR1iu9ISF1K+dTipHO+RpchpiBIl3sT+foKlM1teywG9NoFLs9oSfvRr
dH9fC5M70/RZBrqQ60SAi5b+qnoZYMoS+9MuoZIyNVvQMjnBQ1mG3htHyfdJ91LUM2FKhY2MmlAr
PxocnWUbVcawijzTsPSUdFMpF1bhZuGWZUNii+JEubZOCILckIxOpULkXpxm7zd1ZE2co3n+DhxJ
G2gn3dPEkuGNMz3g0mL61zKHPUXMMs9/G3Pi8WRA14cOxtQPhuqadz14k6yWy+W25GiTgSZ4Scbc
6uYmfiuJbyuTZNML3h9R7rD/Na3Smxxz/IQKUQ75owFC1np7+wTtQ0UyytWOSiFpOTtZ/6E2zQLq
5FD1j6Hlck2vs1eUo3rk6ccSOXvo76Pt3vo1pOCIP/8JmCShi67oy2LcCJA3Qez4N+mTeYZCWNqg
3X3E74Yubw4nUho+m4smDXRQnxWG0v5NVQ1UXccKLW+ZPy9cbA+FCi1o3/HfUlIESgoYgJFsBixs
XmeFdkYbvDiaR64zjZVCi1YrlI0lgM2Rdi9xJbkOqH7qIJ+kzUNbaus2QQreFXnE8CD4XbL7ZNfO
feBpjsk+obvmPRsPuK+bU4w8RQlBSbjp5V3eju59H0atNvYCA75zdoaAOWtk+xN97BRljEZJTcaT
lAQWH6IKxLVHX5DLIrKmo0XrzGrEX5vg3r+xvv3eDR7EQp8DEmsuG1DanogreuGwNkKgGRP1rT9e
gl1l9R0YpJB8ktUBcQFAtKi46A5PGpfNOPrH7Z7CPfzY6df6e4g/JXenTNkg50s4uDNb3F5YVZQZ
qL742Vr5HHIO3dKFlV7atPwY9mj61/waiuL/K1AIXxXXFNxviLUzpNKihn6Yw4sgv8gBopJx8bhL
y5w7NvdMGrH3KmQBr1cKnECDisFdfvr8MKFHjuLKD3QItfZvr9VeftBcFmtPrLQ6jVHbhQ2wWowV
Tl6RB/N0yL24Jx5bt+JduSyAkas2HcLUWuCc/on9Xw0KD9kK2ilVn3LM+MVydEp/nFDz029mRLIq
PouVKCAwvMuNIAo1VkvAgWxg7jz6NJGnoEyzgFUn/Lnsk+IYJmYxODOeYOcz1ZdlY0M4k7nP3OeE
67t/VCpAdEW6RnmYyWcBpf3rmg2bWQq45ltojf90DP3q0L7ayUdCinnrcYSW3k1YbgQPuHwYI7Jf
TRyXGL5+8GliNhSudvqmTeBiyLmDxs5KrloA6wNcatzYT8/5cIfgN+SlUWUk++DXkY5YVsvBxRNY
4RriahsBQZzH6ztcyGXdmSVNa7qdRkcO5Ji/JCN6SYnk1rca5VyJt2Tpd2J6ZKrbB62lshBhxTgD
WKxrRmH+AESurNpqiTFn/+gitp6TdGlZaZHh9T5s4sS+3fHuj4jR1cMfsZQ2FTNI4m3GKHTI8SSg
3dSSEIm2Y3fdOcdSFPztnYWiIAD7wUpF3K856zPt8bcJ//ukraH/onkgY/gUK662ESRvi5cTkyG1
IkgMnd6sVoMlHmSKntj1BCa78q2As6lONdHlmI+52sgKLN/B46f0nIiZHKuHWrJOmaT6cxu4+wK0
M25I3K1qJxSQtfoqBHc8nbA6w4M3erbfjBICG8OkDMVGyAbAFCFGn626o5iiFG/A5D+NbIwf/A6h
9c8/aaSEtRtJtNXBNz38BEOJYv4EbOh6YaVnao6elyTw6lJ5uQQ/ONtYKfMKqNt2TmPxo8dY/dxB
bwNGqvCsNtJL90OJZ1qxiDyG7wVfWb+WcHFeQBmm4Gt5IRRQDbMKDhjG1owlyVxJXFKUc69DX+RX
mwX9/L1hH40UeaIQA8c43vR0HGqijcfAfCn68YzotR3ebIirQEt2v7QNuPa/10IXcPE9J+hlWBSC
mW65rU66eDJix8souaqhNd62FRUb+YTTlMPRr6Y15K7uF5B92a0tyyv3UjfSrdIRRc91mm/BcLaz
MbxkkB7uaKtdRQtA6tuHSQ7bN2uqhP260R4qpoLTQByh6TlYuswLt74FvdA73LNiu1tRdSSenv6L
G0B6Sj/Yi8XaujRtnxCXEYEU0rf71ANPuthVlOonKPIWJH7+DzOfqnOr+rYuBUY/kMY4YMWXUzwk
c3lxlzLC4qU6O5tHRvsRh3oFGWco1zoLzxN4MLB+CZjWd+7KgAcC0uryJGoo4hjkJlNYaRphElWv
nw05LV91YaNIvYU3EvDu+izxPaKV+p8c+A4eZCuQqIw1MuSexNbexTbYOXHEN8/sQ27Zj04r7KZK
05d8ITqUuYiJi0/jYyyahi1u2KpOwt3f5XWLSycaCs9GRpYxfy4r/pLcxFZdbdTNeAE0rsqT0XxW
vEwbT2u6zVaNyF4P00DYgr4pCcu08u1j0WQzgrCG3u+nzXEL1HTgnZSAxxnGkZSXGJRA+zoS38Ir
pRGX97i4NqEI8RAPqIE8Ux5OK45sYW6FSg1FJScKF4rYUJmjiP04p5ydpi9cKVZ5JIoswUefinaG
FPHJsEVYjqxiG4hSarmuFFXdypPpu+mj2WhhpDkbnlArJvkdov5fFcuCx9bpF9CE3ZTbJhG2t+hG
910dzfjmvIDEIjXktECYQiYeW1ISwBIrYu0+1+qpX+9hdZzdwpzgi2wVu2VCMOCvf8caZ0Yrc5f3
NFfnD49nLuHQwrtjpli369V4RRy862q2RZztDDWj3yZ7YLIiQ7Xez0J6eeBSkPHcf4ubbOqkuliE
ROkw3ZAVx/d7HTQmp9bYBZn0vlzSTq6YDYyI4uaV6ciJSZN103zpYmPJawSUHCEY4+IS5q8ClB5s
aCp5FRogNXnvLWbWyObiYV47fZQpA04+txgsZCXxTHC+aPxhRYUn8ULmPaBa5mt7sFUkFmUbecaa
DuJRUzl11QC3TtfUxOqQsS5N5sml6u4+BhEk9x2aBMyMLLwf58Kua1gzS59ES3oYZ4ZUeI30qYf+
AZ0fY48zlCCrhLZ8DR8e1MEOmGsnDqxciydzCCjB575LQPaAOUx+g3Xy76leYG+Z8tDrmIRSH1ZW
k+562OTRNpUdih5WUuekdWLC4yNLkIvnC8EHAfyD+P02Fxfph2bgJ3/1XDklTN4SpoptWN3uuPHw
MJcpEmsyHnHqPGew0rk1gR/LPFGRPhKFJA1vK8vHpRR0xKckJx1dHBhuSClj7/rDi4IdgVsyV5oG
FbZ8Jg8rqHxdGOHVLbP2h2gAn1YVcrZPh5LytFH0yBXdwwG51WI+UsAtRT2pwJ0g+zBvgnnjlw30
2/Kbu/6qAWAZFeVxP9qTaN852ts9jEb7nA4Wp2vKgys6nl3WcURhNYOq+QnPj4D6gETJ/yzWJNml
ETuYEGVJ44Ftwkt04ldBf3vXmT8Jc72VY2KS/xbZKUbAslZ5i5bZzGscczUADKOhAv5+l4FYDtr/
zAZvrc4hBQCukBMJ7aKGsIX3v86tio2dkOxSvH3uGv3lKBm5rcE4vvdpacoX6QZmf4tRdi21/vw4
DfMf4RgGQXo1Tjc31ocCGgSe89+XekNVp0qFET/ge9x7ixq853CtGBTLfg0gngHi8tME4iTYjIml
H40p2EubbTXw3XiAMISkQBdPKj+BvuxzmgTSY1rNv3enHpdEpHwSJQAbLD4tg9US289i3+oBwikD
oeOq+wNyLvTxP49XLLgSz3jqH8RIOSVa+i0x+gI2JC7AEiQbcz9SUVoeAy+yMvunLzn8VkQ58kK/
9xXwQRQLs7swf5WuA5psXczbKGlq9+fVEquuJ/1o8udswGJgDM0Ojl7zdm9DiXeVCXLZ38/4OduT
iT1Zwe14vUa3w0TClkLp3ph8BMUEw5a48rG2JAV2ET/PACdkjI8fY8YRWEkdCFDqWGcVt//HDWog
LGUaMkM/nTX80ZO2XHzd0JMYhXfQrxVCKawG4yfoT51nTXx542vh30bygBsa+gucmfnPpIC283KE
wfomr8CNNlvEvNuZNaE2N1pay3lCLpy1En8VLM7BXPOSV7r1q2W8/qeQ0Qzyy63kNStZjIxmT+Xv
wVh6yqq+m81vJgcp9WjRDc3U/clmmQBUaC7/KZrzlqCFrsjmaCkk9rwU8bsZUTNK5vtznbl5EB7G
YNjoTx7Y9ZsorCsHWU9H594HBL/nytICO7L+nK+8GeALFbCNSBheR8OMYLwRr9VH14WIGQttHPFM
AQol5FBs0ibgJxAK4nKexZgWXZ4eTXhHsGXBu9qEfVk8cNAHftqhE7m0X2YcIXagGHKcqmHanPGC
tsupE2jIe/xtOqYaBskULX/8Kpu7SL+zGKmk4M49tNb37fETgw3T389cHhufIOEAppnrF5hQnwIE
yXwxRmlL2Z2tPlz4hfsZR+HwVDsTwqOz7sh9kUri79JZCyNgD1LcSiVXJ/bxj6VkXNbpKMdv5oAq
4xtyjGgN1s6ZBluQuGHkK0+5orfcIssBGWwD5SHdrpfPu5pwFQCFFZ4SdDlWpqjdl0RtyxoAPV7q
CpdMJvAoVfrgB64pid1S75gh3E4W4/Q1Qbt18vddDt5hCLrfC/tOxeWr93CzFxH0kBnpxw9Mcr5l
Nt0fKwO6HuN5TKzNa7jFOq+mNX5a7w8qOoL43jhu2T2vib1jL+lsZ2cQJqmYpstZlqvxGZQES8mf
XogrYSX8LNxLaNyB4PyHsQA0cY0Y5M11sVHHBBPWL8/IbypHwewhYlf7fee25/jaIKNOUgDyeIFs
wFH7vsRGlxjI9ClPFieYvU/MzaxXP+Kl0XKy6JopoDrisayNAk8In/85D141oHZHFX2YcLb+YB13
I90HDAdLI9K0PrxPz08j/plzJI4BVucLCthm+8VBdXsOKEbtWOe4ZZrUcQ1QU3cT1ObpmYwIgZek
lUu6ySnfW4RA1SCeH8NwPC4zczBmKw/xOBW97r1MRwUMPSorNClixg00Le2DxfVx64w+CYgixUzZ
NGUKfn3njde/v4ZANpzUViwyyP60ptJP0/JOUuqsJbUzKnrlIvWC/4TYtiV63R+XlbbeVa3UAYoc
qlJnzrlJVUBIel2Z6QsN1ZRzwzVvSFog5LNPxXi8IhMMMiiqjfxmfJXZNk9ptJiwC9FSiiDl+iNH
vv+SF81EfPILRV1Iuql+L99vHhvp06L70t8eLipuwfVSxn2o4hJUNCO6dJzxg8Of8STleXcxxBlL
lyiA8I8BPT164E1LizozU14jplPOV+YcXWqcyMePea4TCD1/Wle0EetmEqXMOVUuS6w7WyiYsZK1
SBq5WuaYtyuM0ddqEyb5uJlZotW3yS6Edw+ILtlXJaa7ZVTX+uomXIac9R/oHvBKBZDHtC8UhYZS
xvNGdu4/Hzqijc+PaXAy0RCqAk8FH8Ik3WnmyvHRc7CpMyR82wsCwyGBkrShAFVdtEQcJiTm5d77
uLp5VLbdfRhCsiK6R3ZhUnwpt5g86ByVFcb5GYb6m6jSxOvfIi5udi19jek6dmNEQkzVkCiLCIb3
mvpC0JUMuql8SQKsZci5GTP/aoSp6NPGi5tpeOt61hg69RRN1/swnIvups+f1DERZbyrTxu7zDXl
kdlS1VjhtUDYOK/oCX9SwbweGu+Mrunx7ZgCwGKvW2hLwIrnT8E6l2dCrC+3Bp1dqBMbur9rcf9S
lri38v6x09+zCzdQFMiJP9bJ5cjjv1apabiYuADRtPahuusG6biXptcQHiW5YBHCTZ//AJ3GsTr5
Q4gi6RuvLKCPTOTvYx7LpzBNLPgjenru5VFTe5xmS6y30rMyH056uakwoEOsNTu6B7s/rW37URA9
uVEMp+vEOcZODO0QvOz/lf8GTBZ9/cG2CJZ6AgWtwTUlziPdH59xq1m/dRQXrT6oWf3LsEqJBVKF
snzxsAEaj0G0QRemTSYqGJ2mgDauvVPe2QfkyY80NIrq0HCWdWRtmNz3Cf6odwsG5jHadvNBkMF2
YOgOCVBIyFDPgLKr7zeMk7r9+GeWEJwHxuPQwYi8hRv3R3601UMWGUfUrBw2hv5k6Egb7FJ19YAd
WafsSElZ6oz1gFWcQIKUkeAVlmM8K2nRclcSu64eYEPsmUaA2dY9UaeaOZ09Q7aI+wqd+T/eExJV
cA0cmpIAmq52+JlJyvciD5+065hDYNJIJcF3l1dkSiQ3LcuUQCRf34QvRQejXbKHru/UN1MqLHr6
Snbd9RN9zSG2Qg/T8zpqYl61VjoC3pbgV7Tc4XG0nF+b8dD0YbuLVjjqOKi1KbkpkU/h3YKzj/BQ
zs7sVpU5z12PtyXo/2chP6fye5Fk9ay8s3B55rqaJTW5HdHVRpC+RlVw03aeK9mf1KNMyh11k8xd
2W6D7N5Nlc5sM+7UQdDMDBbE70m1wGC4WtQuXF6DbKCZWrsdOXnbjvmjh/yRdiOo5JkA21B2q8em
Guk5QOwe0qTAYsmt+hECbco49pFCEdgkdaxut1jAD2LGCIYCKy7oQdTXbFHTqjKV1tIzmEZA9Xdw
UGvB2ZE+C/QdBWlN20N0aN7RaafrJx0VTF9Y6MDlUAm23DcJrBDAiCEo8nNG7uWTiieggJql4PA3
096b1t9t9rOOfyfJyrCIOCwDPVIzwGqT1CKvjwDmMJKzUptALXWdu3yAVfnjdJ1dD7r+wnsHi+d/
UNT6WxqUA08ukeU7DPL7JLBvCV3Q0c/g6w5KRVtD8zWtWnby+hEJnb6lbYw3VAWVe20b7c+kiq0K
jc1OOuqfCztVMNXlOlUZwjsDZmJYyklMfutWHBcEOubqx4f1PlcJBcpd4t6Wzn7dNsSBCjiUfD1r
zMwFzxwVgBhX7Ku++z06r3JLDVTPbAY32MC0xvYuChYwydmm9aJ1WN225L0K6fmt7nwPaPLuRZ2d
Fd3Zr+Ng4y308UwPjKQKXynU6EiykH8ApWn2KbPUEAzSOXRBpiw1yu1NOHL1DneR98C36TineSIp
WC7MZhm/gyirSo2zc8Xss7VH27XtrX4PIsc14VFwg213wCEJs3ghU94SJrzNqr410VHo4TINFTkq
FvuUW62qu5+lCOeRTzWwwnSQuXiOP9RGMbMYInBG5UtGsqwWmujrhD6BzRAaurVw+MMYXzkrXL4L
+7IRZUuneAJ8RL2dSRE9342vIU4tc8az8hziAhSx2/KHneQS1Gy8C84HC/iGK8O30L/9hDgkLlRK
azRET10a97F/CE1D543vfu+o1F2got7w7knJ3TVT30mwic+1+8NUxz6jOzQNj4xuUJ/E4eoqjwYy
6auQM9ZICmyHxT19GiUOLUYrJtka9lkaH7BmUDo/wh8SIqZtlxTi2i8aLHEf9pSKBbplKN8EJj1u
GkwxaD/DEbmiC58dU4DZ9yd77qqJDz0wscWYZK/YO/Cn8VEi7fDD0RcmXecy3hyluEA0/ci9XzCS
Eu4iF8sJyzhX68asL9wEmUDP22X+NynlWzNSfCtKcJPge157I9Jp8Sa8ErRKHWAB3MdH+K6qDmUT
6ZWrqpyfk0JLpxKSshpo5cIUF5NfK09ufjtf0B9nLfHszk0cbFa8REhX4fc4GFu9nT4YLxSnqQaX
UdGXD3skMWyNIPd8qhDQQSC1MjmfYn3uWO1S6hRF5E2tE75TU9AZBPIXkK7n4DsmlDllzuK1X7Z9
Pl4OS+E+GrWIUEF7SaUwAY+M56aMHA3Gp1ft3IRzB9ZXmZo9LjlEdUz9KapApjZvbZup7zZh0mAe
+T5hG4SDu17Eg/i6BPCpYF/G0YQjsUFS5zGskUMSmbaYz0KhelyTw9O2tnSXfJZKhmd+w9iJ5dvP
g40MZ1CxqyoGusDbrDC/pVexfdrMu6+k0vTd2OoqsqSJFTXWS/R2HDYaraYH5ualtMjKTSr1I4vF
y2Z1GAD2j6zl2Hthyct+pzAw2Pnb6ZYJ0P9kwmsC0w6Qi1MiV5Nu9JO8L/5j7LxNDAri2S+P4G6Y
8BJebbXpwk3+jtxFbmnm9pK17kLZ2lPjSxf8UfomOUppL80RnAo12jXeS1qvt84SiW2p41ar5hEk
+b4P2b7vMtsyvTNlwzj3Gj/d+7SzY5Xh20h+EcCwwdPgQuUBMoopvlJJTRsUQjNPcKAlaFlUpobI
Z7XOXiYzXnkXubvK+O7hMFAgWpIXB09Uq/JwEUtQ6a7VQgYLnOcGkoduvsAW4VvtLq4SCLhDn564
xBDeZPJEewvOUET7Cs98wFVlCePCq9TcRTD7hYD59HxHk4s5CtUEIn11Pq9l4NyyXPXM7FT9VRdo
NR2oooWk2ShzE3W5gk7LRbpqqiKZ6ZSRsf1IsoMwqur2Y39sMIrjnB1nxEHe8O9SVVC70tJ0bmu6
0PghZ8dr+KaohJeNOTL67IAyQHVz517+bj3ro8zRC7wV7blWCBTXRCvTGL//qZIXeRdZAiR2+I8x
vJn/CrBI686JJ0kLmygTesN/OB19KzQVygbWDaV4WzlWVAA20zcEGsBVGWu/TUDvyIKc27aKNwYc
OhcetDnL/T2B7RiUT01kSMY5YYsS5PQ4Ishpmkw1g4v396tq4Fx2lw+76rZ9P+CjN8h31HdvOT1+
KLkCxxRS311OduogqsWyQLR1jZo3FD7oWhsDJ/D46Xpely8mfdAE2EE2lSXyh+PjQZt1biysJO62
08S8SF6Q7+zU1Ze0Sx5Qjl7LOSOjfHXOBIVKk3820x6OLxHNMxbak/gecw0WHcCw/5te5fKCxfKP
x8plcJLM7nBGOVBi5BtaExjlQCEQNT1OPjeuCdeU05/Klu57PTUhpVT5cPQWNwmrCIQVZJI0KaBH
wDqUmUUGthka3MdPeacdgFA61tjcShO/ULnc36FEsBmJcM2c3ZCwQA7gVQAMoMh7cwmgTkzrDDfK
DFqRk5dLnAFt834wqWxDVuMekDoUtBJBhWftbcW68LLyGmbSK0A2ib+VExod10CUHm7uDMVZAxBe
tCLJ4cN7hHdNqAeAvqY9FPPc34mCRqNLAHe/FiA0RyL6qLiDZCP6h/x10GHE0oDeViCEcohOl3YZ
XaiW9qVjqWjnY2EuRnmtPMe7K7vIe/LGrq1rKYcUHoQyBzoKmg9lvTZwq/pkhzaKjH/eTQBBEjrH
r/WeAYS82Zal+zoD0o5rXGzCy3T+Jpzazfl7Ik3RySWtzoGbZlxKWcrRnVSfjw/XH/Tbh0zBp7/S
4qsbZR9cv3JK02VgGNaVfwRL6GoTGIhLB2XyX4Ph5arXjDmrLO6gAuaIkjCGQkmE1iTumUOqn5Qh
OWU841RkRllP9Vzc3XqNmyt7ze8Iz9/mjHxUGZYqClC2fB2/QTv5C11Evc8tPMKECKw7nx7X9VCc
yQDckBTjF2I7bOp/sVV3GwoYX5RPxPYQGz8nfWVSkUPop54WWHt5+ha3ajE1YuZ0lsx7FJyV0oiB
3hCOrnS4LreMw6hOahRyJx09Q8H3dZ/PTdXiqzchnGEVXOQZZbVTAxxmGpsjqtBvD7q/Dwl4SVXT
eKmuO9z7G/vyNnwcr00/fhlJrS0J3OTPC66QSOEORV2Gclun4fmrDegr02OyLjvwRGAkOy3evjXK
JxkR01kZRX1KZpe1j7/AKSVlcFbTHMCNCmTsU1eJe8Pwpay0T4h2QAs2+qGinHIZM+oGNoh+O3CJ
hEQBRPnEhgN6yJhsTgD2RKvqBltMDydHiRT2IDZ1Sj302TKgtYQ04on7fe+TanczJvrjF6uu77h1
PMIdo4TIpynJJ0D1h7clrZ0X1pdXHuDwoquxUn/grx4Vk2hh7gsL8dItHkcVj7yGQa2jvn39CTmu
aeXMRQOm5v+O9+77g7nfRm+MWJchq9eziOU6GWdJ8BWZsNfqghmnwu9tnl1xWsyOs2fq1TQoC8Ox
Xb4ddhSRxWeT9A6Hx3UH3u8bdaDZcN4NnETLO8ZG6ntj/s8NbwioUMqqNVfAm2ZABvNrXdpg+ZXm
Id3jeWhv/VZyPH6GzyoxC7lAXbabvxrIffKF/53ooY6tbc8us3/3b2gQ87YtLyVo0vOB/zZvXk3N
FcLr1IEztfKrCYX6ifyxJC8lyWF0B2BCUGp12DI04acmBkArGrU3AYO/7WdD5M+EEfaT+erX1J7q
DXMrJO1qtl5wXRki6thXm4EB/Bo29mPy5OgJVDrfHQfJretxRQmqSZ2YyHSgDZFrWZq0DrpfWZPo
8K9bftNEBVKiC1Ao8ynj+DA8l9rr+x3xSgN5vjdGyNN8ubKx1x3rd8Bjoxjo43C+0wKP8OtyqI+1
5o1WBWOG46yAcdXI7pakiBC+HTMGMCtI9YyV5n0okq5Lix18F/PEXxZqGfSEg9WKrF9rOn+P0MsX
F9VR6eREOPtNGYbQZihAVzFkGyzl6Ou42xEgoy50UKlUR5pbX1ivZn/LXsuAUKDV10HDKLeqH0Km
eLBj6i1EMWguyReWcpDdQYYjlK+CDBJyosgfzCWXrRW3Iu0kJzn8udStCUlT7prW7q1iM08mXiSt
Nb//oH0oBu0N6iQCnqe66G3dOfAG1xyKTP96LfqCD+5RzKopLXNl1H4RHWGDmltNm45qx0Piz19A
zgeCTlguXlP11tMADCQ8AxjiZ3WaKVUR7/f93bhjdtKhSq3qMxbWwhNVuBrtnP0I/G26fDXFyQKU
UMoFDtS+hF2gS0N7YhIkaPCBVV2w6QOJYpBJ8mAg8qEO3wAgZw2AyJKiPtG5LR910Au7fkmL+tGS
EW2BjHf//GxFHUoe0LXtUfznjFaPFUmJLAKwrgV6cw7cXzz2Y1QBYQfCzfs5byvlx0hDmMhrhdyf
v8ZV7u/cm4pLLBN488Y2YlLVSgSIb6ON80LF8Rm8TWDeNLkBoZIiSsY03xtOKJL8kT9XTQf4ohOK
Y7lPOlL6beEpHScwJbtPEU0aeA9PeZCavstLmeplheSh0dirIcCRdHv51s8ZyUAqUtA9ebdlk4vx
tquB74mZyIEwvJAyPzaV2sIQtQl8qBZxgKf7tfkEPkNT73Zj7/DxfNnoEzw8ImGQsFT/zNdFscwW
+Hdqrx1ngBTvr5ZFasfcDcSyzusfP/NJ/d8ZYxyoCgmNsqPyljH173Hgoi1R6XYvY8+OyxiIqVkY
0/8/FBVyLFjeilNd+0TCV+qII/I1ZsNMgZwYzfGZYtnLTeXws7MqOW2XPULoNHOKD+zaUofVVCHe
FC/kC5UDCBjrUmjE/+pn9SJ6zTTT12K2brtgz2HEkTRpfbbZVkG9sYePggyetVSZJDmEtLm0lb1r
oWH9gAlh4fw7KSOgcKnwPQXrtKVcBGvKJ//di1PScDPrQA+mYCbYeC0UFKlbtD2n/ABAyHZeHQgW
Y7oHLh7FPDTQtCicsiPU2U/yVjSZBSR7engEmdXQC2sLZQNQFAPPHI9f2e2OsMaCDHG9wC4YseIh
iPYBhAN+mrwP5YRm1WvWIkttmDFaNjbhlQoRzxtiK714IxgolySSekQ1OcFJLdJB3uyapiz3hEM6
Z6HnY0ebGmLBbFkrc7mCIKoWPMy2ANzoung5BgVQmJmPTfzGr2LTLSQW+TqyJ5ymPq9qd3eQO3XY
6A1zDUY7TyxIDidwbgwwy+WZVmGXdaQPM1qeF2WoynVRzCWDSxqAOmjDGqtnC14o4ZXy//dJ0RXb
kdzK3wROhkRtn8zM3I/lf6OWmJvXbipmtzlp49I4dFMKRH6VBc8z1iQU5tlGI6o8UJwG4wlyViWi
AAwhxZgTxpBkdRMHaS27wXkZw3l5te7bOavVB+WD6SGcgQcW2EReWNnliTwUk2XiBnWbWrZ/HAPf
0Zo4FFZaIgPJItzCuDmxEmSpUtmSymUiy3heK60zvy+cvQhMgvI9DqTMUFaEneXpDkuN8V4Bqxu7
eQeGVc/70xKbuP0cb8hkCielKzTVvrjz8u5dqgxRILA/9N1cE2vifCynGwtUBuFAk3gaGxB6BrzG
8fDlbx5TYKczSsHXPA3YFYk/dFWgD3hbdKtLZsAbYH4GnBKDjQKV9PUwU3ZUHX3U2BqL+PoNDGwA
Ar0XhK2kqWM7HM5MJy0f/HEpq5xSuNT/7fvVq1g74aT6uUGLc8sqV6Z0L7ng7Lw+1SpNt1MuEeYC
Wr6NPb7tgF0Q47RoxjLhAFBz6GS3fKoh2wYFr0sGcxX5jOF/mOH1mfazuMuFhn7AFJi6EWDbfMDO
6M7t0IHLEjG+hiblJGLvJ9za4EUiBFd1voGF/M6iNFU+srMV4uxtAKf2t92pX0mT0qwxyOkKJtbU
oCbxLhtpTpHBWEZZy/nlJdhcMJ5EbE9WRfx4dWpNULD5+1OL72qdZFMUHfhg2dzS6f0y2Hy8Z0e+
KaRLGfDIh9yQP9FBiXLDlvh8oYNaWGwQiAn4DCqu9clX7kdSXDmOdO7EZdDFbQW/oarqRL0BEsdl
Lqyy7iIYGlfSP91Tisp+tNyp0oIpLorhJfR9olQ5dpulzXGrMK7QidrtRyaOVlAAq8Fr+6mCLzax
LQIRU0skXSwC/qUvvfAzSARWSakGq1Vh7VlpB8C5LLP4pT8XNUXCFPOBkFStOxZn2oy9ZANGhjHM
Mc36CX0pwVdq1eehncXtlZxArX6eutoZjLiPRbwKnvwZcx3pRXFcu4nTLmHEvVWhRdvoP4us+mwB
393pqClL3Y0WTmDXDe61Ri1YAWUMK1VAJjntJIDlC9foturCMLuB4EscKeIu4zWYPsI+LuQe5zct
cL3AhfkNuaxVI/ykdAFKK2nqiwmzK+/8qJ0/kxctxLOlUIAQBdQWumvtp7ooavt+MYN+s4UT68N4
cAW36ppg8WKw6DdFjRNdV32Odi6msvtPETQx61wgmtJw57LewTzKcFTxCbblM6psFUarT4sxxO7f
EiPkirF+UaIwhN8NOzwvRCvoUWX317G1ZwqLNtKOv1AoWaWMccMNqwXJiTnLV6573mF7MId7a4Ix
3zgCPY8A/ukhkPIZmo8Bvcdx46y1prAOHFz1ulByxFHuEEFDjwKZ58EcMQQY+gaPKEVk/4LfHzFQ
cRAs7qlWq+o4gghlbD+0+EKmcFl0BOnUqw5v8u3zjRcEplF04HfX7PX9Q1sle90XQURvogBKkd2A
OdWRiPPctQPBwj++TUHzb7vO/BiLZfUxKC5I1m14kB6/rpcd+wm/w1B8eUgkCYiajMx3CFs3P+qK
upHVKekbdndJJvP6tUUdASB7Eh6Ocyh77Pjhpj3eS75avDvtt1z+Q1zNje/IjmIANOt4XFUz/1WA
3gW47sufrBaE2KYAg4FazPa/Gl4LiK9CBqeHvVjIONoxAovEwDRrS2c1io4+HAHvPi4ePDob5dIr
bxf3WySeNnYn+Vu3TGxvdsgOjCtg68Pxzncu2hQhDx4s8p2H9Afhm7YJc5mxctHQEe/+EHQ+PcsF
equKVbPI+HCrs2KpWjN8XsyORGUDOdj9DiT/9bM+nJCK7T5fITDTkCM4ETEBGzzcl8K6KMA5QvjS
JoucruZNeAx2aYE9jLR8OUew59B+CvWbnXkPWRwoWq74AViEeDO8lzv20eIPbjHg2i748R2Jk2gi
BimyjkqqzZlJ0fJ8N9yLBjHGpJFcxsUK/NztP6sft1iKelY0S3refIgtXB7j9blTYD9l35KhUqX5
6xDMI+Juusj6NBbebP5F+YkxEvH6NcezzLf/X0kqPnKTP0vFOGd3SsYSrO8TSF/QmvJ3lHN4gwbm
XgW594V/F9rXODfZFId43IeokTS8e14y5Qf7S9v2fZoiduQkABdIrfdyWWeZgHUl+AQqn+uSG0y2
++zYI4AOIlX0WrFUxfyMnORnNLa4dFkH3T1mhiT7ksZOZtEFfT7c4kJsTEDXF9tZTxnSXVzpPyz9
kjxKd4BxFxDtiz2DWTl5r75+905vLWrQpnjOcatYbEwbcmm0z0LeyDGCKC/jZyyleu4FaFrrUMwA
rM1NgxWC7zhnv0mJp0j1HiRYp2cz6KjF0LYRo4j0LOvGasRWDtIDGRRZe9X3I8sJhiAFYxQ1s71P
E9AsPCzX81RaaNua01Y4weQuSrN5rTYwBecwGy6XRWx12uyVvzs+fmXlbuEU06PgMc20mnsvXx+7
J5ucihctHj6sLspiaCEqjc+fZbGSp5otBhbj584dR/Cb3M47TdY7onKG1a4BKVI5ErT0gE5wIoe/
Igc3BJ+sHx2Q3snzeN+B6ELHA21Ootiv9AmwApZd8wGrF/8efTy0zpepmfI/obZ3G+gtBea4gBi7
nY2VutZMvhw46z+JKY4D5wSIwkwp8lxdkK8TizsiohxVPnv7HELMri8S8IOftMgxBhEkkrx992Xa
3K1v/Sxgg8jwAkNQePrgWjxUtjoYXxmSzah4wFH3buWhTVlOKeKlW6CxlHEvE3exQvcwB/C9UU0m
5CBMJmEbqhE5DyaNrI6UCgYjjP2WKQi5cLWKnV7kTdIoylF6Ko9JxPRC5bY4h8HfZ4IhQ2uUGGcl
UX5q0Ks45ENWiBhpVpjo7ZUoTZImqMC3tZ6PSfojiug9HfmMBlgWf58m8Bne92qUcNLrlkpZJc4h
dDR9ExgiyHyEAkUlw0zWTLqnVyXalGi3df7xaU/T674bny1956ZjRdeFIauhKQVoXeTnGEGVWA/y
do7u1+C0m/OuVvMjA38h/tGbioqBfGJdKrJdR9BLR1sthLgBpvgD68TS5vYxE+rPBG5MR4slSXIO
voXDKi8nwYwF191DrnzpQRt2Mau8QyglftTVuFeNUIwvWo41RwOxaOUwQBfpVi9hMMfvE7/V9063
SCuAgru/MuhL4ytbe8TV52fh1fjgLiJAZ5FwvXSQWOxD1LWRZhw24vu8Pe7B3rkcCKRGFWjJiTKA
tNVpNtRGtPAeHpQAy0bCxJ63xyqA+H7NBHQpjkcQcQnd4wWJvztMnYKj4mJ91w0JcPYHTiwI4t32
B0oC0dExkRK9x3pAkh55z6CuxS4mzU2lXxZvRXfsL4lOdn8229/oBlOO1Vju+gjlDvWFdN3XqYyt
t8qH/VH/yzmihx2dvwLMLSy4GmNfLvQUq7DLToN/BVfTpc61sPDw/q0KvfLSfOjWvE+TqZzFXAmL
OWpphQQHPHPZCH399/ue+9fttxj+cpThL/qi5Pb9EcQvDvF0o7brjY2rE0UeKFaPk0DvZ7tm7Tj8
ndIVgoEmRSVMDKWdG85er3lVfaW17HQAEUX4+Nw71a2+Bkn235XAPEx9Y5fAAKM6IBBqLqWzFFTv
8ISIgksHOS83wg2ymSpoc6O8YP0PfnPf/+tupbI0p7CYVO5ZW0MPX03B/d/A6SkfZrnfXxDpuEd0
vCBD7zFNLX2cgOf5j14P/dgUG0YisWxk5NTQopGSxsIyJ0jVPIbzwgWxgEVcoJjBaxTbMCNJ4g3z
UmSYz3PxJaxGeHKufGYSJSG+IkopiLq7zIQCbHblS8Cmld/ATOrl0CLzoHzURCRdzOsElTzikLG1
iVpaWhmRQqA06lrI741+gYJdJETn8xdVJtd8DRSfYzn+iRVmPeE1xNZsnTXhvF0f1mKjM2fvoUdi
2Gw7u4KMk7er7lqn8sfPBFKZBB56BO3pP3BHg2Xt1h4mM6bRLmdsTbmIyXZoCZKSi1ljW7D/F74p
E7gMK0HHpglp4uHvePq/tl3oozhTvXQ1LWlZ6rXDtnCnKxjiLNUb8XyIvwnOuLcJUotBAIBr52Ud
UW40Yzhs/WCRdN4GX74FAEjbyXwldIY5Mq9PKmn8IZMtqgOhzHqz2B3X6xffMIEmerrXAa/8ioTT
GPJAYBjP3pFYyBPHli1+JvyvGybdWb0TyAcqHtLWvG9jecFAIpOzY8teVR6lIRvhduPbrWwOTTJR
54ujmVSqXHBOFDnscRVIf2aQRz2+dJiM5bEpfL+NgQ+fEyIY+FqwhK8DlolzWGt2Mo7KF7VlfiU3
R326/Pkrwme53z0h+7VvAu6X3iotoDJ2F0eR+eLkNgZPkja9PqdG0Zt0/fs/recEnIuq5fk3P02b
sO9RYZJeNMnQdyNilvSLcnLufEzPQywxNwdwaQLMhyMejoaV691cEJA8nbW512urxJUEjtPjr2X0
z9WUIwvyITvOzvFRX8tfJNhnasyj03pjsJyhOrFoxl/PfMUgvNhXxMAI73KPvTxgULFzp+jw2a21
Q4VngOs9UQ1UUozGjFykY1lSWUjWVCP0N/QKRbtoLmjbbXJDPRAb8RJlNEPV8OOjDymWlr/6D/f9
uZC8G0Y7v/0SmBmM7v74Z6cvb0ENXy5lVTEslOAvA+HjmOVFPjk0Hs0UCT1kbSKzGkuBj6Uw8QH9
OP3Gmi5omlsywO/nGuYOqY8iUaMybBJg9tLRGU24WdDYqmYfkil3CN3RkMwB9ygRWnAqwZPp2r3t
XBXR5lYkow9lAEsjJPpc/FB0y0w0PWtR0n12crg2e7EnzC6TvuaP4t+bt9J1FLCSRtRKXIoEr+3Y
71x5A80UPws8fa1dpVjP8nDdf5kZ8xDrvg3sBaogznPyJEoOegxloCCp/GrgPgtZ5mEEoTkwgKFa
Nkrd5l0h3MZz+yevbKN9cjL7wVv1P5XgSLqBhZWjnRnkwc77ivMirIoLMwkXVe/f6O8AmrytKr6e
ypfiWQH7GxGMNG7IH7Lfn/szVMq0NGrETqfYDsUTm8b23VL/gKng5gdB0mYvm64/n4J+HNxoI0Z4
+vvqwx8ZjVKK+SGvD7h1JmM2ytd3P9XOXnnuJFOf9BO6TIU5YWWwKLsHzN4D4f4rM3OoxupqhxLi
YcAbLZXWuVXvZdt/EZHHn0T05akRnXc5CsAK5FsAv+LodDRiBLlzz+FKaP+8Mj61n1hVHegfYGGN
HuN7CZ6XjQyf6Odk9J6ieaWKhb2QLNQASP2guyMqib7IGFXCkWPFUZ6ABZfHuS+ib6K+c9lOqhgd
EckZ6I2aWFq3G7WpYfAuNbDpHzeqKWAvfmadmtRzKXLV/MtwZ29QngpszyFsDqeexk7Gqov0ODDG
UtoryIFv8BUzveHtfenpz6aO4q9jALKWevU3nrFc7vXQaAAxJkXuW8aVJqXXEQrIhRMKSg8M8nb4
HKUWhDc9lQ4fkr0+eMV8eTUjC+t+UmDoE1S1rGM6cIWqk5YmQOX70DWGOu4rKs4QSYUcdZgux6NR
p9lWvZOu4uCGeb2yc3An5CEVxpTJCCxNDyTPtQpBSf0Re0Xr1ZQlQbKT7SD5raMqNPyssq3zr+GY
+RTp+80vemqipRUP4jzXeYVA9d8JCO47ML1WmBWl/z8/oe6FaLUJDu8V/5OuVza2176Is4hK1P5c
eqQGAwyEKvgk1Rimoq0fk+7QlK8/1c22kNttsXOgGgwraoX46igKl7VsZy9QP9l8pPQJyP+CfKZz
KzZISAtu9+c7qCdTzV+fIWVg62ZJ8nbVXG+RGaJ3Cgnfvi3rGtkMvQYQ0iCnYKe6mBKZkpfA1H1l
9UJNgW9BkaSRPYJCfBoJ8QlcnqmOrMYsGAptzvuG82xYdn0pXkw32lNi9haCDYaUblF9/uuKHvhv
rswv4Yd9VobYlqp9gDv29OMBoRztEO11j65exjc0uQzVD6fmvAIQojasp0XV2+Adoemaf9svny1i
wzOKGeTS7teXCsrrZdWq/VGY2Cx05VHpnGTlidOf96UNSLPLuSn17Haj44C373Dl8t6n/mLk9xbY
TCuvsi9DPsydVypoi/gW3f28OWiwL419BDlCziPmlgTOGkwP0TsUOBsX+9Akgyvz8F4IZQNu8D5u
OEyaevMe0wjIrqqLmFL1Z5Br4PTAvmWuIM2KZyj+S02U5xuCT+pMbDtN3PYU6QOYkItvOx8K8xRE
s1FtW/DHQzF40DzxERRB+cKr/Lb67TrnSE9Stj+lpkzVzAKMkpYcLYpPVVHD5pycgzKuE2q5JAQ4
ACWbNrr8d42oZxobafoJDPoY4gNwU7Hxfj+jULY1ZuwiFmdN8ZFq2wLFrB0JU6cjaowZNBykNGTL
Or+BIqA2hRjliePLQ6Y/TPMcKByuBYiWkL896jocKyZqDM5KNhipO4R+b5UmEJS65RwOw1vmHRiw
D+cOMEPGlGhOWfGweoH+03xEKGqwT0zW81D2TdW6NhNmYufEGMErtscsR7z9uiHYaieiGUxhrSnt
AXo7WRjQSNBxk/4vIJhLi1Uni9Y/y2dqY63IvuXvIcTpARLv6yzN0PKD3KbHMWjwc6GIpgSxcG6k
NOjXvoyuwawrRYJ2ity0jp0JduKYFVm5S0FClACF5sTp+7jd9rNvgWrXKEG0OgiGjQOxCwVTcAq4
ZH+7tAkeMPO6gOJpJuoFs/5GLIlQTu2Pc/0eRJHw/50ACd2CHX+e/C4HpfQTl4n1gr1o5Vlx8zOI
sag/YpCJTdjntLzqS5B5tgTclcyDmt/y4LJSlK9Ta33rqUqHCVn5SoVIe8VUvIouDwYbfIThJZt2
U39XrBnunQ3uSZGNmy5X+e90W52XoYRllCMqnxK8Fiee9mYBpORIa/PpUtERbS+n07r4Q9xxz9Qh
1zQlQZbdYrywkzbWrAkUTrq055UPjra/5JUV+3tWCdU+1G+zszEelivJOrFANDZ3Ea5XdbMtYt/v
pCHGbZD4qXYmXqCCKLmk/TD73C4PSrbK8yYTYcaDpq5YcQklINJPXl/OmKiuYv1KbLV6B3mj1eKg
cPcHu2oiILc9cYHrvH2H8CziyEOMMeFq+DzCV/P6sxi7JXiiUYBFevRCVczozxerY9fVt8zFjrX9
k16Faro1V/+AGJE1xdG6nE399oo3+63lG28H1zhFqrWpVHQsNKg7RCC9xKKRNphUkrq/99H+xOOj
NwgbJznypoKBwWMXvO3XzW6ZSP14MxyZJqUlivPsSFrGNSzcRjmqz8eTfaWgcs2urnz5a1tLyluH
AB/niGJL3nAnP/LMv9rYqil8V5LsOXj0qxhmAHvXMLSbHgvwp2S8jV4kgDw0Bxh0MN7SeGM8RKf3
Ig4M0FyL5TMCdvsqH4PyyLeApv6fah4OkDua1HNZk3Q6dDU4gQxoGqIWvDkzeDLNXHXb7mtpfvki
xR3k1dieyX7cD43hadO5f3vD681RX9gWRTZ/e9bjmIIzJ8/YQvsmsswcxLPv305KbJ8CZznSBReH
m/SU8tJEI1xIOKHi9/Wono7k7KaIT4QhpsyHOGynhUVmFfQKSW/fuuT365QhqnaN7rgDfGXeDsk9
KzKbv/L+y+fCWUkmVgW2Vv9xoE0HwYUUgCleXxJeIcBIy5N5eRihcpXNGQFbxY0TAnUY02fFhWe1
cXqZYg0gomm2REhg4u+12boDHipA6UHohC1wN2apOf8aqhYfNFgSHZ2lMkBo4mp7hu54qlWDRguE
NhpLfng4b4FXVn4m0VegcoCaEuMSQi3lwK57B3+G/YR+qjOWqimXZqY3BmAe8KVvxiH1rVNEK8oQ
3qP7hnOFAHiJWPqWKfupvnQaTzr6ad9TSiFjFRQkSLN1E6ouxIlOwfSa9r2RF9mZDNzJF0bgojGz
hOhgnElTh34YOCUE/smT0xTLykKVmqbiLLapK2JCngK+SIWKHJFMStfmPbMJ2sqvy3r/KOCX0gVC
NhuhBe+Mc+bF6qH9U+6H5I/eiLU8xLqSZMq/wMdWh0otMb+C0FwwzTn7vS2nLtPlCYsyVpjSiaS8
lHSZs9PzIqeOKosUdQM6BF4/hkDLUXvIxeHBwW8h7leQJfXnDZzZ37HOfDCwMqOYqcYW/KcARVny
D59Tcj18CD2A4Wv1SLKo7PQ5Yy//QBVrxzojNWbjIOTzrAySDJO49oqQxufiZpiW4nRf5EjtowNy
viHyUlxcfViythjAM7hPHOGVbIXuPVDQpV2wiQMp+CC37Qf1B8gYIyXnJFpTZI/9+YUC0ItNT03K
S2IzKExaXHoq/zwGoKNlu4oWbxtkJNsh2F2G41pbKeITZQ2E+saM2x+5AbvuuTw8uW4xkQm7uHkX
5hgyoYWepQeUvS9ar4GVsZvfG/qiaBfaoTRlpQxTkJy2xPXzJBx1pE9NW/G3au/KCZgZAF+Qy2FZ
bMYtxP2cxfS3GJJu9sUMeQ5D0JU9D8xi4yBcDkxcn6GpDMjVmCwNm4KxeihsJhex5O5+QQ1/6Rz6
PwwH2jcufdNdw6Sehha9DP9IMvSP+3Wdy55BGYHWdVCPlSMKtasMrdaKev9JVzuvwHownE5cNkp/
3rypusd+X4ZvaidEeuaJnxXkcBC03Hrl5JvrS0+mbbVJxJZcj0CQ2FVyHDcCG0cUxrvcsbPr2/Rk
8IFGsAuwpwQ20mCKKldiQ1ekNlu3Qy3hWIrCNJl7UdzHnxX2KI2jCc6oWnevcaTcJZShAZzK9WDZ
QdgPHK5nDPlhg5aqnPTOnJWrAEF2CxQMRYmQerEwBpRCQy6a6Ickt3fNqioJQv7M9Zscy2LWPaaQ
mn3qSKIFztrh1ddK7m+TRJr5iPTdqJRQM4Iq0bCKOxthUsGvPPMAtZCXfkSNoKJwYDF1EWMDxjkK
7yMVHVQDHibrap6LnS1huoTgMevJP6wEZb0bx2IfFLNGysi08DI/fBESXl4TW4zojQVmHURosy54
wd60yyAVOdnq/4EAVU2aj+cED1JbGem6PMe8sSUb/nApo9OpmrDpSpt7H3DFVCNkZuXgGusvbbsD
sLlHyq438bz8aT6vLuhRJusECc4r+T4KGv1bPOYHWxUl5Xzj48+pCaoDKRku2MkBuC+koIfKdlJ6
KXyo1DgFhpwmXgrfD3CaabOMIAcjTwRR4GoYpuIG+2EhvSjKErcsWXYm5dcgOQSksMOg+gCV4Rr+
aWPCNwdsZhCiV4XlOGyAn/4yLvl1UZ8SYPLI04GBbdT3FVBZik88KfUCq0OIeuHMzS4k8DQUVdPl
Q+QaT2CHEb2wq+dhepzy4Aa5xyc96nWc8DghHwYCwPEmeJ2te04srqWkwSwoiw7J7G0W2AII3AEG
3CRdQqdwbbIaS2yXJbC5fAYu67SZe9YGh/c/qT01i2dGdIrZ8qSPlKQynQC2FRJJBq+vk0wGT4vt
gI69TaVs1v773utAgfsc6uFERH8zyf8t1GCRxLObFQwF1bvGSQIvbSCCDT8/0Sfl+PJtdWkVei3M
X4IJ56aA7WjOmd0jQ+6YO4lACjGiamL3cnSvxW00L8izsArIBUWlJQRpISpAAreXAzNdw4qzeSs0
ezfc/N+iuxJdYpFR3YmPUgI54+NEUQNUumy/1EunqMLOCfna3sIYy/IL9ywylOfTta3K5NUkU643
tvSlsvmxI/hI64UvLmFY5RWWIbDqQDDDJwZlcN3bQyxJgrYSe6lFed5PoWPIfoBWv+dRRBOMHgcR
gawTQzG8i8suBvZ4Te6aa/XWvHMVC21GZn8qYefpB/fUUR8vKOjqpOo1wP8jUFz7DanGfWa7rXGb
HqAtNnWndD4IovbizscRblvWa8DPqMPkaxkksoNMOm1PwaKtwwxRzja37BpvHOlOvgXaVt3fgyus
S5criafWuuPauyoLx9kAFfFRVyYH3Rm8wpfRb2zZyxzdyelZw8l/pDCIMH6gumc0VF9oXGZXYDoq
palpEz5gjJN4sioU9ckd0ANoB8L1tZQZD36aSzWmmxawePFEWbObkFgRU2+HN8NsqLOho2VkWjWG
8+ze0amACde2519Kmu4vf4lnTWawtDeMMiue0iRohrD+nLOtA9tt7QDLMYFOc6nf6oGHnIA3cPoe
/XNdNbZBaEjYvPLaGyUdF9AXkbLW773omRg+aqE/iPsK12LvG1tA2BVDUrfIs5lwpXRQygWLKj01
Be5af2DwPNq2ysqRHAEOR2tgNAqysDiZUDM3d5Xo8qDci3/E3GDVeh6gHLaO4iuIdDSJiib7DlIF
TSWh5NxX1kGCyGubkatDZz9d4lmI6fovCtBp1+fxGkcOOBzDYqctubcFCxI+KYbAK4puiCHxuOBi
wl2KfpjdNUs9AOajJQoL+s74SzA6uDpObNE7oWRDFtqGEM7NoN0/QADlXKnlTyMFLGzW9+D5g4yc
4gXe9Z7NWhfE5ui031LP+lME+iklqps2FoBTN5F64kpjid+TW97BE1H3WcTscxLTiNBZudtD1wYO
vQZ5sCdq9qlB71B4K0xcx5SliYoNy8lHbFUQB2zDz+5uDhW48M2HxuZkRUVGpfz/2ExAc8yDj4Po
QRNMPAONSFZ3eh+NzB9zWF1hMImSR1o+14k8F2DyMHw1WEkNvpCwYj0NyHNQuTfOXlLAn3ygKzcM
MBlO9UGcGBtYKKhs3MSSi59bQ5FwH+3bOxvE21GI5xotPIW/FvTouV8SjlZEA80PoOEtpMU85kfn
a7PMYo3MC4+/dD/iJd0f5eBIVTvXnopg/qoDD7q0rNQrduvn9GqQkREvyOH9FDNzcXLGxLKKB8MZ
7eHctG9fhSPCM8MpaWBOi3vHRm9pNmU0tjQRshx46PSPRbdA7AI5V5fs79v3T6SGeNuhiHMZ+rYF
encQBI11mNf3TSkKycTnI22rce38IT7rVahcgsEC/4E+DgSEGHnSI2Ve3nvxTJSNfFwC9ZeoOt5R
o5hsXaP2pd4dRGaW8mSy/QUfqoY705o6bcvjRZBXXHzLL+mXUwHMJwmHvVJupgnpU7oXPWFZgRCT
ZRQ8ZP6To9McdaoyM/aAC8F8l4VvRsodqn/58wPzT/HzMFy4LqjJ9JhCrZ6LyCa/XydVV1NCObKh
Ynws0BKV7WXIW0ez/6Lo+G1O6FDa6QQWWznxSTQfNglhGaCDqLZL36HC2S0ybpLiSWaUJHkwAosq
igA1PF5aAaFQZ/FX4zI8oKNkjaiZ4VCWroiSdrzEaB/I7wo3LBaVI5IYMiq0i2JBoVgaZKHO7Z9Y
dh5hBs3Rn5+w+w5yxeuvlwqXJlwemuUa3Cry6QZnxYDkq7WmJCryN6Mvi4u9fZmGrDukh4ahqATN
Zhn8KEjatgMclSOaEg4Bj9KeytxVVfbfGkTf2hDgDYEXorp3Xlm/ADtSUpryrcF3vijWUub68Fln
vk2F1nMFUoownum3RD7bHYcTOAC004Nh3cJw62akbC1BeYfWBcZYLT/8Q4Y3kl9JgPo9N2KDHXE4
ZRJzor5HIyQaH2kxHO80qzNpd4BTwR6BAeoOQIfAqxcXbcAMbR6m4WpSHiYUbYfLmPDwSTt9hv62
zqltIyDydifakGZw5moXYxpxn2E7RugN71211Gac4nWLiCmk2xNTeJibkmkPT2FSC3gmL6LdVERE
L0hg4D8+9sR6vMXofh8Zg7gwhXZ9PODNUAMj430soY5wWAgG4WO+fNMz9qKiNOpdP368jCErR6/p
/RL7ixTUBVurCHB71eb4ie/WoLE4pWEuztr01FSZB7hx+DiAphm54RLAjs2IKfMrkvl+HQch7qYD
AL8ym+4FuIDUYVX8WgqV9MsXzrHtemcpMzBGSAyZNsoG0F3Z7Rqwya87n7ReLbNbpOS9JBY/V7l6
sPx4PHnQcz1fSeUxJ3H+GdOllxQVHmYcYWsZzwd06O2USLvmCxcEEL4db9an40uJAmU7gWdysiHx
sendAuHSfPTVxKKX8cBOoDLJgZxYDoAhaRs+INiuAk+nvWOJZt1Kf1ZmWY6YFPUUGVh9p3c8Momb
YGjdHIvG5DwOWzslZkKXRO4Qi+WqakVWKj8e3gePXX9UzrwT4wuGN3+auvysZkJGbOc5h/aod9hw
xNdCvIzGyFCn5jYAX7++4zBUxfWaC5T1dbd3EJr5z8o62dvxWWDUUVn+290DkTXgGabu4xQ9HZIB
D+6iLVi8O9zTEao9Odp2Myk2iavO55y8XBKkWiOtwFPlz1QX9EwvTAfw35Ip6bdVHdZKH+MLmsdo
lalmaW67ltgIU2P/aE4u3sd6P+ZDIDY1IW0JRUnxoSAp3crh4cYbTrrO+rrrff3FuM/yXQyZXIJg
eC/vEvUD0Up34/rZdEKvIOhLIk6EebLXlu/hLZAbMmUMpv1Orh1ri1IwGzofcIGT8hOr9QPBxvUM
0PAhJWAy0Ba5vIPsAxfiRqCO4eGL1X4QBfOgs3OPIeusUmFYZmnb4ceKbsbj7NV9t80PFubWiBV6
vq69sApS9CvHqRRJvxBGkc5+mvNnBeCJ/t2XyDD3XcyHumUmaiHOsCzglhZN+3+FtzkXU93s1//S
n9TJ92EatnyIw0a1G0zOjrxnxQhi1o4fzNL/pCgWtPOlhVmnh5jzI2xcmasegbO2ZmWxVFZD83ja
aDZ5LNTz2AGCmnl9j73NKlQiLYEFUbvOIsPKKc5/OJ0sLCFpBwU1MUGu8IbBZPvc7DjoWjJ2VVbQ
4NhQbqIB/eh0oKz/WyxiGND5nuZwaaGjoyAlm+j/35T6W3dZy6hfKQ+OoDhadkPmuCBAjjD9ht9n
MoN7/6iDE4PGrzriqXuxXXjLJUD7im1T4xa3uMZtVnQFMz7q1sKDh1rL/l4ep+u2hbBmfZqdsMhB
gHvxMsldA1u131Z9H6po1Zaoxz+yy3iV0+OKRphGwLBzct2JdKVpTVaZNjZAWxJ51s3zIFeDKAnE
QFy24TWEcuvB/vTXQOKayVKDVuLEdgyNZOrBpDEHgp5t/aTtw5x7ASTskVa9RPVVxbPqRG5wNB0I
e6jv6JByfvXoXpoB59XbCLFP3EcX83PDODak4quhwTtqrnb2cusxjTUgf2eka9fvhQITZ1b0LF+s
WgaSoArNUYvIw/wPYfwcWzXE3P30HaHaWbQMfnQLQkBeEyGsICX4Y/Vk3MTz4lY+O+iIglYaOLp8
cLuque5+5ZvIHIii8jcZnweFDoood5bUjDpymj14uui+n00W6IPObksBGdsFdtDLlA2zhpsTO7wu
ZTIL5edpGMjjlZcALH2X4+erUr4ONhWcYd1AugJvNuwFIUOvUGrLJvFbz29oMrAtDzi5FuOTo476
4ec8GkJkykzet2kgcqtcPzEiajU8S14jkYwkoLD5JfeUWsV3kq8Joo76KeMQ5MsLBzUK4yQAkbGT
0+Quc9jmkAikcG6z73dG+NpanmDf3XyH1DBgldFRfCrMcSUB80nFf5aYr6I9GsizSQwyosdusp6X
n+RFFgJxDp1lhcciXdKWVmMEHf9I+7qqNN1bPe2BGZvpGjcP9/OQP9+I5hEZWbM7evVsUmv1UkBS
VlrYvIKCI/5aKQhF2weCf2b2OEglzDdoROTwiTvdY3DS3uF65A876oS0fu7vkQpeMFJGzYSgwwSj
3FfwJUyou2RG1UjOt49n2bfwn8vcLOzFG+wXZ8hq5hsPgWHrKaAKlVq8fyHlUn4EFOEsUDugCxv3
hwhpyL34dfw646D5+Qk5LLZwkHdGLrY01axf44YrXHQin77yFJKamRI8sFWGbP64uCq2u7D4Vo1R
2bTlMXl1iERbBtqJxi4a60LliJI7hEPiV0KA8yrZlVaoFnzmuAafvTHAMMx50QI0UTnH5SfFwOMS
mwa+ViYc2CPSv+OCZYb0jvpCUg85skZLfMzXoqTS0vfmdCqDJIcTMXlUI7Lr3SX97wPQlo1mGEfk
iL/JGNHga7ZnnqK561NRzkuYbpjAtvCnnX6yxZdXbuvxHvpTiPtaOVOqXjtjr0HWtXX6ofP+Sjmd
9v4aTmsPzbGPK+BaPisA528qn7vlrk/YVwpBjq7lMOMTPnz5Lp2OwRG2LvHF31g3LgxHMJ+LHVuy
z+NYIVFnJIli8wcvUGczjT9OC9cHgd+EPz5N61B87NWbScbt+Lak5scFx/nVEuFgp/iGgRmgChqu
GHoYUTg/ph/Q+CCTTRwyu+QlcOOQSRvDXPpFrIypR4bgdULwyAOZ6aPcmkktDtK4MPN7S5/v70uF
5ydt6vCHMWuzFESoRXEREWtF9jvLUiEXtd6eAeF0LWW2tb7i6Tm6n9Pq9zVtsAsYdHpkqY/Nqoja
FHhYtjituMNUl7hp9zf0mIKmXTPfnWnpBWLb63KYglcFLTCghjrMmD8pZFkDdN6DOGDM++OgHOkF
eYEnX+pCgv3Zx2Sre4dcxLEFsCYcaDnAHuwHzLf2ZqPhm9srRoYTeW0BJEaWnbxXkZZ0ZA6egyrv
L+d3ITYq6mopLNEbubepQEoDuPM1/JBo1n0k+EdHbjfIlOneSAuWHesyyKko852fzPxycBGkBtsI
COrr43n110PPPxD176SfW1BJcvY/okp+EqI7pS2ZkLj7+h4iikim7X3l0Q2/22l78uI0qGoOggLO
VZfjsGePG3mVM5+MIi37qdlNWE/avyq7d4BCKix7nALHwvFrQgVfskIp8wJbRlmPeGWL7sKiPbCn
Lvo8oll4Df2wSjtOhdYDDsuwv/sh3cBVdqQUwz8eoyHjPddKChS3d6eQ7dsAMPdMvYDnEZ4DzHbB
jHXz42lbfO5n/XyvE22ZH09oHKMi/gkCO3kM3uy13ZAHikkCq1dWrcT4aIlPJYxZ/9et3T94hcYZ
J13k683XLBoJEWw9LinKBdYjUX/NLAsggVdx263+VUq8BcBoGDx2jyCrhDR5LtpV2DLIb54av/pR
eoXWul64ODV6C84+uIPWyTKcbqsPcXpfjs9WeqfDMUTU5bGBOawcCCq+ACljRlh/0uGAMxYGN6OQ
ti335iQRgBd2cwxTe580zvwgqqz11DTRLoCe0vzXjYQWQBv6yWCx4xCvVzJfrCnjTjoquqMLOWUb
bg6+An1f/xvCSEVQZt0Q5hqCGP0c+eEGVyNCAV4/NOt4rfxUXzzOCpNiDKCYvOtSnZletT1mI2KR
R0cO6vMNo0xBEbgR+ztF2OjbbZ3GD/uLYkhQChOOGnI1WJIUYoIgzFh4CNAWIH4ct3c7kThntRom
7UL703bcqqNHgsPtkucwT8+58wZ9exq2rpqpIh0juG5vtupoEjhe2KDUF8g/uuVfRX1BUq0JzC63
vtbjErfFgBzhACsml1ItYV1LkcckePslxHDRSfEDICEtQgo0ntY+JVAuH4CznGofilN1EMh8D1Zs
ZriYuBD6ANnEQY0G05lF4XzuoCpoTiZ0P/yzmvsMuWaCWqe3nWI2pxUSNK5D16lqbpwf8/RBrTig
Uu5i0WdxPN0INdnHggm0CKshqpQDEX9ZoDU8GW6HzPrwrP8N2alRiFgkKjH3O7MpcP1DnZI5Jmdq
+EWNZ2qO65VHVC6WP3/lat7MO/qiEpLzfBO9ZnXf5YVbHyFKwLkFScuzqvzOHlyic0kyxuac5i8x
M/RzWw9EKcV+6zSwK6Ef2c6cwbd/PU9lvUROZmw3Aw7/+TEnK63EcOq4m/kChwELBMu7IjBQSRsx
tox0smmogKwpd+1crfP++C5VReLmY4iv8+9moKUbjUn9SgbZxq+tmdG2hqr5s+T2cYHHZryI0W0D
bZEgZO57EsRtkr+QdO4sty24W7wSfs6pYlAAGU740h8SS1gEaOWkCpyckBfwjMvVSg2llHOfXFwN
Eo00kdxy5pwqcnkkCm5DDu3pqVgrNb6YyU3a76fiR/S02ZHRB+igcHo9yZkgPbdZlyp2nl5q322Z
r/zCMR8r7yk/xdN67pNKtAcXaQD2TVxJ6pvtcAiLCyPfGO/nnC7ysBOvypuIFSwdy9405GyUBAd6
rWAYIfRjJCTY9i7b0NaCX8Xs9iwSaHEOzu/5RKZmMUXQCQH2HK9jbebZpZGT1NHk6g3aZVYWPAb4
3fK6hURka4EA456OJU0vZL8jrya4pjI6C81PSePWe68h5m8LLGA9Pm1+Ou7tKGkYCKvrYqKfo1Go
XpLBiah3m4IN87fGcPTzWoWPbykTom5wUc/j44lIDR9BmLUVRZQioG+PIaEinEsaIGVQVEVQFE2L
pHJWKFvMXATFqbiWCCiD50VwIwRKhSY7ulcvLQQVssWDzhS+UuCvlSwCTH4+K3obHHeQA2RQwTSD
gjZkXeGyrqjFHe+eAR/AFZjbrSzmEXIHQrOTrBeDH/6EGXcYW9yYnaNSp9rqVoJ9b06RoDtTF8ck
4ZXTVdIERcUajlB2IQ9spMLeqjJpZv+J+ZGWKfccPKvvTANGTVuGhjbdYgyiKHxTl2yoXiQMuw90
N7E9f3kbWlkWtwevs200ThCPGybJLlikfT0DOMf/Td4lwdVCekrHkuYihuCVS8LwUgP21jLNuSjr
a+Wq8Eqp38XkM2MJoAG+Ewf94cegNB8tGufke4zdUR9PJS9CuZ3zQShrKp4e75hkAlZJ3uxcgzhD
Db8KS0MGUF7DS73nS+9D30GEYKyne1n9qiBT0WzWn/jAzjNjqbVFBIRudLWPYajFIIYHm3Kwbjhv
qEE1Ie9SzFNty3TL+mpDuJsK6cvbKw5e0abZwT+3uSm+V/CDc2og1VQL+Oo21tZTIiXbSbH13HLS
7uo/LiGaXTHPA7Gp57UA/ZYbUI7djqTNhKZAWesYfcdbPn1IjgfUOKD3buRL4AAyRhn2wapHwb4I
IBS78TAQPl/nxZoKa82Go/gG4LU6XWG3/5VweAovKn9f2gPHtC2JoYUmkgTVVZI8bEuD3mUNqD20
QnHFG44ICEPTCzQUYte+90wKcMgqVYo9bMM7YG7EwTZ3t7fVCFvkYTwN7DzZlmJJbmig/KM5oze2
cZ9rxbVVSc+jq/skbgQEZvs6RKD7DzEvrrgWLudb5ErvQuJ1qU5eusOpA8JMeZbaTNTPdoEbzh7b
nYTH03eXFUI/pjh0BQCQpKVpnCTYTzwJjcgHg32/vBtpTcIJhW1frgxBx3nv1bUvRVsapErWPtKU
fr5p19SLFxeXOuEuqGaGkzdzZUv6cdLOSxznpgNZzczZGJ0EI7kwKxmvHFHRk0wjD5srXWjABA0u
E7tNqlN6ZHTeJ2AGcGnBWdg8Inl7Hv5uZHNpiVHgStsWRjToO1pjPdAFDiQH+U0t4GcC7DWOluHJ
Hpgxv31TghzJZB8+M//hDcxizadwn2aS+KYC1uvSqgzMjI1EZP+3h7EeaX1xn2DPCgF6j52vmvq2
lSNes+7yAMc7NCk7TwvuIJsX9s6s7LBl5Wey73CioylitpOOlaI8E1uXp/vW/XPyvI2Q455rvfqv
rpPuy/2YbxIR9iPNIEmwvFD+CXepgeqn+RGArtnioQML57UPBql1hJa2w0UiJ8N/VT+5wf9u+Ui1
f/I/h4iqqPzu4h629q9FMrZjzNZUusXWTKNkeia/AsYkwk0/lF3+qmJCO7CXExyet15f0VUfDpgt
3gtF8HhMsulV3MKP14o5hkzRLtB+HhjpcHx+UHPAye6sUUFzm1n5kZN9jO2F50tfmThVWfYfyN6Q
Z+cJUOWpWpcldGejJtLJpKV48wVz1m+ijUO7qu2NAAQtpIRpXlnBtXASJon/4Yazok+SOM7OsVpr
+DGXjv82tCf4M/w1a09sBKH8m5s9BiaHbWEtm+VTWofQzPkHxcv1K6g0piCDRq3WaGq19uZ0pYC/
vDmsJdsumGw=
`protect end_protected
