-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IW00npK+ev8YWjB1l1PVDJTpVoEK4ZLcIabHCWDRcSr7GEmj7y/Uk4Bar57HUD4OgajG84Vssnkx
nYoe8qjIr5ec4h0vX1gfIwZXf0ePORYWGQoIIrFMowqyZDj3kEpWfSvKliq2/x51gHXwMNZKFAQm
On15uViyQD1ye/s1AWlNLPXmthXbnARa4tZeUA4W/QaqszFN5SJFoj6ljW3yz3Oss7KylWE29ATR
Rs3gVwvCGtT+Dwf5f3ZW234PhBQSrxOIR/IsxIgnu/C3OuQqZxeqIteldqYFswX1pmIWRTK/nGL7
sh+Jo8NjMDeB6Ysw0Dn65PiJok6wWcYafMV4HQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
5+vTHxc6BLgv8MjPhvq7ACmQboyG8VRU/ubr5ws8zJZRcfa6myb2ngGJjzg/PbZ61PY8n38NvDQz
MrRwNU+3FctgxzJXCiRN8JjOCceOGq6m7wJozfOxUo/Dy6LVsJZCC7sYg6WlwdRt/tea7ZfbbeN7
kraYjmAk8pUmhlmmAYDr4cSwpmyjymdBHh9D5YwQP+kMHrXGX1M8i3LTOvdv1Ttp6S15rKIqeClJ
yARggD/f8pvw7cy1C7n2Zfow+0b3TLf9F/Yo9Zyq/XWw6mtWvMKbiUR/DU/oc5Hw+xZcD3Dghoh0
5hM0TZIpKRlDsPgMnOR3kh5sjw9e0kvSSb+tbI6vg8KUADvQYXLmfshLNl8EAgrvMXTOXPIiJcV3
eKQ84X5uvTpUx2QQp1pCdWQwb3GGDUntXn6AoXTG1p9pm+fe6wzCqnkUAMFIx0uQDhfZc9rlHvzw
h9N7VI5pGOvpOZBLVQtIrjCRiA3cWswAU2zCG4bHfvQktRhesN+p6xbX5itpi25tItkQp90xB3RT
0wyJjvI2PkhLZb6fl29QPk9VG1DQn3WnVBZDUa/+ZpUHlhzTnolraNE+leTQIHs+G5VGVDKe5V3s
GBauzc445OSWwK0Ua4gUs30goWt7CZvzkIePQMdX55CuGGnTSpPVKPcY7PbLMuXyGqlZWK/l7zQN
rpLGQjuK5xVHKaKPOExtt9CJgV56OLSgIqDBXWYdP6hW02ZUpES+9x6Fwze6CefiMpXWizDcya1R
FtqEXxCeKRwmxsaLN8nxi7BjALZunHur+ls7r4QVGAJHzo1meKm4QEHRl2v05necYJECopZQ3m47
xZ1N4SbLTB39w3/BdcPLU37Gf2Mf5jorT/wLj+IKpe7aHv+rW1kEgtinJYszh+6oNbv7co7GqnlG
kYqup/Su4JK3+GftGJmI/+4/QMUcIZ4iFnTmctUTo1b/8YpSNoVPtTgQdkfTnmwiUniVXeY4h4MQ
9Ae0M1etD7bydMXrDJXfhwhRUhhBu+R/5GOqgXE4IRSp63s9Zy+S17u9OC8+1d8cVVvdOvC+HzQW
xvUE2CdL5db8byagIZaS+vKWaD0KrmOKVxs9c5z3hwVPQ+YhJnAuFmPAbW48OzCn8mynoN274HAa
HS2jHs5djQ+sLe1P718HfsXtb9F4upWbIZRlwj6QaXlvDhtmpR44tjwPrFRB2uQGGnE2RMn8oZet
FQCTV8dLnhcM6lXMLZEqt0KMZ5As5CDN/sptyk+ICwO0ajrh01cIXm/Vn25GiNNn8yYyFVdtYM16
CzaXdzqoIpCgXq6lZfehGsiMeAy8FcKo5W3h0vZ2Bk3L+ZYM4tUC26R5U6wBEgntKh/aFtekiLxw
j3vTw7bt3ldKehS9XL3pg79xbihsYdWsZkkkBtL6+0zGEkBfO4ZM58xbB/oa07X/wGZieFcAXvUT
XtMlTJfOcy9OLcD/A+wNFE2j1RM7ycnTGJOGdcat9rV30PJCMy5Z1DuhAKlx6tqkoZeq9y9Qgski
G9nwPBAoBN0AfwwVcusjhkhQVdZkf4ufj8k3Y/dcVBZHWxaz7fU2sZg2rLd/Wfs82vGEnd6AX8to
fr4Ic5UWKBDkhMr7PyEtY3tVEl0nWEujsKi6a9d18ucrybFFgSzoxqKxzdDqU8tOvRqXCo1Ij5fJ
f/fcZ4OdmaLAFJWS6g8lx+YQ7w560YMsK0iQCZBCKSMZSfuiX6Qk+Btjj2mIptDGLNHUsjyuM1vW
mxJ1Ihbj375p1Z/B+2czckMD2gduUTNlIdZS7N/8FiPVP5sJ+HXbnjazpVFuMt4KMvbilEDSabMl
AxnUCmjaSVG7aJ+TkLheaOdty1P2iibmigecNTssLUyNTxbxygBdfMHAK2rT/Q9dLGj2F0CGzXWx
r0Pg5P4IF1wHzUxBIfEb8hJeXoumGeGvHH5UrZjuVrC9pIN2SBiXFOKhTwKcLjIN0WRvJRJrLRFB
epdmGrllzFg2b1ElqAkX7Llvha+tPjp/YUeeu/ZBIJ2D/hIMqN8icohUu9a/mrzy7izR7yW0H3FE
NF5zB1zAfhI2uE7sedmPLFYgVNchqg8XEEIs63LlC9mWMTEPswmI8cimMS/Qi3z9nGi9FfSTcV0R
tMIv2OqEayQEJqpSgVEcUB4IgDwF7KP6mfBP8GZm9vKJSbCRGNdzC35bPXG74JOoXELJDOO/Q2Hv
rH9Muj9dzwX+Qb2KknWxgRbfaNhriSNIzs6CtiQbIgFEQUqkG6vlGbApnRfsUGHaPK/F5EuSBO49
4nhQMNBGN4huJmBGGEoJwwAuHi+fyNKGdjqmdi3gVMpeIwGGLmx9xiJtvyAYi/7ahrQWxK6j4LdQ
4DbFhtTkCpLMtbxjlGTdWLSlNxZ9mKxqSDcsUocZNY7Xk6rQjBJnyXifoyUIQV28pPgzztI3keh+
rcML58EIh8W+HtAQnuo0CFYvkVvN0q2FvnL+E6JMz5kAaw9BBW3zKnPNzDPQBhJoaHLfK2Lt0KKX
iUzOB/JlcB7HVwwFCR+VgxzFVELrSZIEw2iMHISNFNtT5Y46e8izJV+VF9mijFPM4xPH04S4vlZX
z5csKoIl4GCPdwcLKp7GkDOA6u5q3HPK1g9BZe6pIXSRnrZ2CcL16zTMKPrY+xaomw6zbJz5NdvS
VBgqrA7fVIX8/+TQ6ulYkV+SiStcktdOkpDrnirTAT55ilgY9AE+DWtxKkB7sTLzt7IZo4JVqoIe
/7P+ybSCGIrMZsjP+sNnSZz6xd3mRi70SBKD3yoCj1BUGpOGYfcBpX7nDFja8ayYVY6rIowYiShF
WDj/jvnSIk2CoMKNL/su/M1+j8Z5CW92Ze4dEcdQ1zOx2JYt/75aeQqdwTw/pY29pkyCA6MF7ofo
Lz8QjHXpgvMExiDw6oV77amZdgEXtA/HDIgpqHdu9nBh6gISPIbRG13sMTyuVfv+94J9DNyW41fv
/Q9VpLwXjXEIfXWkDXz7CKiuixpF567lDReTEGQb/lAxD0ag+rygNzVNT8uplRgmKr6MkivW92EJ
4S3/W4njpG/dbNlrTHTapqeu3q+QWZZOJD85JMY/RvYEGziog//IMmKjcUMQxxzmkSKLEE4Bv4l0
WwPyQsi2yLDHk1isppd5TWGgOdQxbjSupajNTBr088XWUpcL4idtyubwR/IoCulETvvff/gCsimL
Ma6t+JV650BmR3yx+kcKHkv7t40GK+E8nvSzT8a56C2vdkShq9V4khkalWQJhIqSoCRG8KBNqVU4
p3sl4JLOAXHOiy3VEgRtZSR9eTe6yONhRYm/OMuvBEWiDXhddc2XdNJ9tWQdZbZXJ9h07YBGmyzx
Ve62738EK7xlu0c1+lQisv2LkzcjYimzsGoARmsrKBXA2iTGfdYJCBU6vPc2WA2YcoYVK+DrOrW5
bow939N9TeXOIh5/2tX4kyJTkSktJpGIBPhssqENgbZm9zu9kUIszdjNNTq9TjibE1AjrFE0fO2p
eXNWRFPwqoYFhBxSj0c8cJBM60Ex5fVsj8xBo3tQ+vGiGgs6rhqLABcoVnyzwayjBci7cLvr0UDY
U0+rOBb3OpPNFKA8LR6x6ThBchw3weEcoZh0gdUP/Uko9ozc6p+d1Bh5/byXMZG88W8ACLLTs8Xa
gj7w8t3z6uK+I8G1lV9kpYnglDeSNuLn/QPPaXpfyJHbc/TYfIxvcgp97LjaL14BM0/eQnMr080Z
B0vD2hrbYgMtrTGtRCuUPnyNZ2sS22SwUjQJ7xcApQaf4wN2TOBn6yInXzrQJ9K+wmjU72fZES5w
si2XCeoadIxXec+MECQWLNicV/lzvYGnHAIZbYv4oliJ83Vrj3o9Iy+Vszuwu9FogrFwX3nJ/9os
Ear+6I61pkcK3noCGQZFb5MnRStje0vqjZkNwWkl32XNEUWcQwVsrtgONH31h7eXbZBs++ioPBtX
mD8EiEBqqRL3v0iaCGcRfyKK6s6y0UFCMSyV1Yqx/v4hsqSOycB6WiXNiPfUQXUVhADGkBfoy6Is
be6GZ/8LWEd9S0A8yeeJQYsvd78LDmgZ1ftfyLdnArO6AqgA1bmhuyftvv/cOEHSzyxMLv6gukm/
P9QGlK66IoRQHvnWjYjsMCzZ2Sq0+H6EyQH2c5WI10hnNOhy+JP4Og5fcSWZG6+WZDtKfh5nnLn5
C5VfM0d90OjVvncVB7fu7z4Zj7HPI0Z5C1hqyzL0U9GWT8ewAbhtLfM/iBzHPJza9ngSz6RKlUWC
crUqzjONHfwoh8vGzYUH2DHOH9UTQuYrHr80U+OCQpzHHQRBvVt/gw4W2zX9EoExSkxdKpYBSZGa
G/qZQ2KwHf647XbleNgO8gwHm9bSb1nQTte/y9j3wtLPOTOHOJ7GGl/SnbvWmF762sCQYZJeoz+F
TZVGxRnd/1SDy08XI2OlgfFY1DuuhG3YNyb0HcxUDxzpVoThy3R1vKh5qzaIYLqDcAnylQ00zUMM
jLj3Gx1wW9VZjFr31qvQK2smkSRBiQZilC5TS9VvQYe0BN28c3RTRBYaO/wcIdG6EMrnfn+B/GoX
7fJWO5bhgGkRQ5JsRNH04H3cjv6Xm6xQ24C3UECtLxrmiOXdjhWl6I/VbuXs3V64thny0BAa/LEG
zymAhqJiYfVbr+ifE5yzAXZpEFx2RkoHLsvCjgis4nMjmvSc5xC+xiUISSgK7V2vldQ9QoMgWU/j
D8vul1ZRh8/I0IfSIv5cRsGMzZLjmD44Om4bng5VTQKBtGTHQEcBdTasEY3D9Q/OC+mcBmBh18kS
//kTxtfaQZkDzabW5F94GCna4XXmU2JPzLNgb3ofEWQCsv3CpW4wfkduDzTwHyYSWY6Y4R/TDf8k
RS+mxGHJkGaged7oNon9tRuoDzoR+8NIJDydx9PL93fMhAK6WbXI4Ghn2m+C71eMLr+mH2NL7/Y6
z/LjnEDzrWt+pEN2ZlsPajKwOCAGvDLGhZfSF30U+K45S/xFg0lKSSl0fStHRUDfOZ7KCLdRevpf
Wtmhex/Gy134BHJoQ6H6vJ64ly+SC3OHyEPgIWsV0CK4/a/yDIKp22HQ+BGhJG0y6ALDO2htT7cG
drpwvMvzfVM2Gr9oSR0T1VLalVYQNI7Ofwrzh1H9lTlrAvxPXaDtL1n/ZSn+WRUykcS/MbACFVr0
jziwdm21BPiDbH7iBJZZpxXqlmo3GtUAbKy+Ybtb5fUPbvQ2PHbmCrEsmersZCH74KcyGV1HEpd8
MuOWUb6F9E+8MDNxbQh+nzXZulnK6yYIN+Op7c3Xl0PJ4wahUXLwfrKVJU/Zi8VCjdVt8S7fP/XO
NImhdMuI1t2hcg58Xi1TbnE+ceznOODpDBYc2NoLEhbbmUVwcOmOqx1h2LBA15yxT/Iz11dfBxxN
5aFroG6eX9chYhJtgDUKZVvs+PFA/bZsqzvKeLjk+nMQfW5BSYkfcMQYyWjuPl1VMXy91LFHI91J
HO08WmSHr9jps1eoTBkBQr5VJBzm8GkUlPoFsm+6baDAznDEAK9Qg2hEcIDy2b3IQGjoJt97IksH
/EocGvz9O5B+/DJqY/iPC9xzI1YyxFn5BNshSMT5dYLj67uNxL8iq9FZ7jeWwlzW71y/TS/WPJaf
SV2ayZrn9/Tdb4xb+Xv1c4RLCs5pdIIybh125r5dceZvlZIopGtvp16ZRFiqObesjFzOwtPxZFGD
GwGuWH+P0RYGVUOMFF2XX4xhg2jYxHY0xbK5ztKoKGhHYlqFvBSBTT73In1RZ8TJfHb4ObM2TNn7
tnFoa7yFCMVhSmyzOJLCV0qLifPQUzJunYlBUS7XN2Ca/QdgQR/EBMzGWPBZkAbo32SYO5dMn6/u
kSOqzCy/uFHbIlAj0XYehLQ1JLye7CTLXJAFJuYmCuZTEOiFgdeAJxDxpjjwMJUQVixnXoBkJ0I5
P0jzBPz+TU1Nn9DgcxOyQngP6eeSIZZ8bY+7fVT1Hs/D64xmOOX0SaH1CqvYu8SaBpq4x5psbt+V
s+gF6npT9UhS+sfJximCyCgUnHmsG7LwaWf2U2Jxa2656WgUS+9I738OJSS7fIt0zrmw1DefvbIy
PEp2Vp+YhOjdeWCyY16WegQdobDXvF9mB0Kk9WU0lr0IXOt5CuIHwCUYUbZQYZUUj7lQFMnnZcYN
gFIUdVSbEtd77m4YD5ubqXzOT5xDrktdjn9gH+pPYS6QFBWbpB3wwNGqZ00LGcCZFtVP//9Q3U4X
TnurRxkoUWNd60RlSp7WMvkNx6LdGQ3/1MmkK1UhEw3vMaBjcbls+r5HwIyVUPXxDKQjw72mueB7
Gox0Ue5AnkefEzsUDZ92CBcquSNIfrVs3+QzVZxtDVApZDS+pnh1iL7KEd0J9mY83Ov7bpoNfNwe
yEyTJQGCJaiAo68AomorR73dKqfVQsOW7UOK3qRjaF3kyZW3nXGSsmkJ3kf/IJEPyO6TgLhV7pOP
0195xmIgtOj4qgoph0De7+r/jXsxMw05FDXuOrw/rit/VF6L8c+e7ANZa8Kvpx0B3n2VltRXo6Yo
cMM0MG3fjNrG1WfvyqJg6EVe6H30sLe1iKL9HceCXqU7/H6ZnNIIeoEgzhXLWwOwcCTLs6lb9eYV
IzXoCfp6CyCs4WNuIK87TYwkqq7xFFcKJmK6fNWNvM6vGMblaEnRDKVYnF6nxAvvaONxfDa/KjUy
88FBlhtmmESBCVS/hRIrEQGKBGPqB/DwAB+c1awLVpxMJdkgKlNekLEzcXf1pK8HmSeGm82+zkZb
szG27d7mInrQjus39yanerLEXrBqP2yT8PjauAc362emoO49Y/Ip5WBTgZaadFTLX+5JXiQUAg6S
ZXVoAkgWqXvjdz4hZBGp7xniDf+0HhckMKzXiPolyPepl4FuzWcOViMgxyB+ee9drSJnXxWUAUKd
P9Qb5d2j95cG468Lwz4TJZcz0ZWziNa/SjFXsw/ZcPbDzfqQYb6CUWZ4XMySIi7hO+7g+DDmlQsf
O1ptRCZVjLEVe0L+YzZCpTKhkEZJkDL+mH3+phNN7RM/HnPLskr+AFqpS8bgTUP/mNhiXk1PRGQ2
ZQ5ZsrKwRw745rmRY/Q6k7o5fQv5A0HmH67IBv34713obdRAoK7CaP6APh2PqhZoE/irV/4PKrlu
tUmlQFsfJ8Wa5bqsEMLcouhz36mBvDz5Z3Mv3D91XuKYdqmrtlVQC4wYAvibL9GJE500OH39kMd/
4Fx54MTeE1zwGzlIFSe6i8TTW6DWerEFjJNxXl/eKgz51dQ6zDwqlS42rTdgrBj9BVpeUq4a+MVW
t4X+5u1xZWa7I0El3EkDX/6Xyt12fwNLDdaicGbOWsyLjpo3ENNRCy9P6Wp8chQemGLjqBquvFlQ
V97nMRfJhw+cTwSckoF2FoQno07F7nAhuUKRYiC2xKlb2WDfbjaFYUhiPeMfGv0WYrrffVpZ3rEs
+AHleE1ueoSmVli+Hi21qT6ZA+LWNwn9urs8y+V5GDd0RrG1RPcH3t1FTQFfPKvs3abFe+XQot3A
OEe89fWPFMTnrT2ebMVDTTw0IqjCjRD7ZAhJtEF9BD2IsFSYpm0wBczaVHNPRhl3mt0gC0eD+dHy
2dVsY71dIPQtdm9U58mMrEgZMvNsUO3Oekx3hvs2srqUwOM8KdpTay+ggjXS4fgRc2jOr6kYwcS1
8lsdn9hR05vWu/XCo2898ZICswEdkoh1iTkuDYDxQQumwfUQ+Za8MwthcLWM5IJ7bbg4X/uDqh3q
bfUAfoIUneFPe/eZf1PRPYegmDXZosG6Yo51VItnT5KjQc+5Q0Cf+sI4lZZN2CrWl44JqdJnen+T
hEIEJUfjhJsTAT38n5HIAmj0GZhJ/8lEJSShkYwOq+h9fh0juiIYcBBE9f5b2tJCLd0qwYjElz2D
/5E8qKrFQP/RqeF66QnMGNI3HLOGGM5xeyPhlf+iWtudl9J5PqpR3xSOqHFvl1nUP/Yd+a1X4V+p
rP1SWrdzjDr8+1XZOrHV3UuDefrP5M1amKHvRehJBAK4Av3idkpBDfrxQEgImKaxOZ+LAzxkSbId
dcATZrrCN7ok/qp916Wzxqkkrman0amfbSXPnubN9t2zfIvXwjEdWW1y8Hr0JkuqhttJuxB5aoZu
2+3+1g4jOEuwNGBjA/Nk7qxf7a8LSQ/u51+sLyGGrR0z/lc4T+DyWy6ajU9a+/hbN3QPckVac0cv
mxk+/wr+nTeTloTVFh4u+mtpNEI4aYKmk9u5rDasW8Bf+JEmRwk8ELClUGkicMeOVijt95gjvXjY
3zxpe1tGLZogysld5afKIzAKkXO2X45NfXtIif7fZNHMmL8pdM/WmqdA1ts0Gcg7WNnTc9Mrg/7m
Eg5GkCiyecubCCHC9vSdvE7emG7+M1jGU3lFJTBLpUUgKJLAcINYLlSuUm4Mx5mmk2YorJl05/u5
A2xKjSpppsuJ81kcjM9s6bRANS3NXQNNdSK+jDN3MdPvN7ABActkXrkQxt8VFB1htEc03yDhmIJH
trgx+u59kRfXRR015RFK1Bvjc0l4gbTQdSdCKvENWE6xOF7GgHBVvE5saMYm83vWG2knRgVSnKgE
jRzXCnupM6lq9ISGWviqjuXNIZIEZZDortOdTcBavr2ICtPjtvDovtec3h07yA9vInAdNbY1ledR
OADRgHz0fvsaoN2txY/yfMRcyNifuE+u6jZO5IboF/C4DJdCBeH+W6RtowcxCGKskyyuleYmRN0B
2Itbq/1hhW9EbY+cWkXAbvvRYT0VVpSbeQVAovgsGfg4IfTyHhs5sQnjA1Gw0bThVAk5Cz+VvSDJ
hdhjhM0LEK/OmKxCUka+4vdSaq6gKxpE0W4TXPmWOqCfoMF7/C0O1UMQ5FqnMYo2MOCIRgv/woVu
sehZiJymbq2fyYGQSVfENLNKhsrYWZD8HwlTA3CQYGD+wjkqpJ/0SPzXQLMFV+1iztEk+c6QHuuI
r02MI9Iaab+Sj0AlFnP2WtRnSkPv/qkpR0RXQzWhLFFmY17TwVMp8PJD62XOIL/7SQ275bX0qsrn
6Hw5LB9zPz2jYVgkToEbDUbrjSmW7vGHAP5jK6iU5BTIAdarRY2MzZ3NzAXHmr9OE3y5XLGOIq0R
zmkXCeACcxfgjwdKCPJLEkmlOu/bnO2QN/2iORHuXMWAH3dhBZg3VDGXaqEilZBJVx5N4fGwZogH
AQzNj0oJkDCdrYBGFSQP1nc8sy24m4PbL0kFkuk39jiuGO6sk8rhQsnEzDL7k2XFLhipJdmLG3zk
FaZeLEWludv1NDtKHJVwAOuixpPSoKAe20oIwez6Z/sdvx6+tNmVx00hMvqvujO/RZGyRKe66nNm
VWxNEbGgHKBd28ZrWdWXqJaFKGfc2DVBtciSYGPsAvrnBuZ+ZPVcsYc+t/nPeEmzhkiXkCsMPExB
vk16Ibkuvn9/UT/u2PgyFOhPnc+XOBr3kps3AsbVw3uiUMVgiZ5PkmUwFjl8SLFUTNlB/S07PrVG
8WUXBiJRCS3O6aNGu7pwtneCbkWduFNKch6m2J0Of1IuSPcrAwABVBxEuxH1Uzc9xo1IUbgdQIeN
pTtFoV6EtV++p6oGnvWhBCUFb/KyulWLtSupfvLQgxUMUjzHnGF7ozGkRhikZARbL3tBX39XFdQ2
NiVgtzMI9qvs4uuVOSxqooL8FNVx8S1w18LyMTzm6AtCnP3Ac229wE4UpUY3DYU9YVZxXuI6hA1y
2uJexuDo6Azo4A6UPadVagV60OVNwZ4zKSGQL0U8MacJTr2e18MYV6GAIUDI15ob5Cee5Y69yRFy
WNFZGfwxu/vywdDeE5SARht5MowVf2juzd6PnW6XRpz4CWmRDliDuwmnSA3RRa3youB8qEAUGQzM
jUl/XfuuevX1AwYj1n1olNDGFTjfvzTr1IHiwWpKIEHL60xxzWy1lZw3szUt8xUl5D0bsNxTzykN
1sLr4/bAH71gOmR/PnwNSOmOYjVl65xgyVuArvE6qcRBtjKhFbHEBeBqNne1oqpGjvbxHb2pjHFF
uyF/bBpeWaHr3kAuZ3vGKYqGsz3Y8/uZG0WyVWN3NXsdUlDR2trGgZHzWIQqFVqUIbSllaM/IRH9
K2PyzKflyOlMMWlAC/sEt3yasaqNtduwXlEPLD9hWZTQPtYghWe6A+rKAlzAMEEYyLJ6Zhh64L8t
cnQbQnT8Pq8IwWgWkIY0B2xa3eDOtaShSBSHqelAue11tQXl8dHgtvsO4tGf1bJ6ig5Hl4wqfSsD
l+pC5Jyzr8ui5fE+epUHfB05NdgmEtupFSVvCosfKqwOH2eaYKPl5sXopO5kfF6U4fFvn9nbhNzU
LCC+kVAEAdlIHgvCVvJGNh+buAZQXgjjnIlWODwJl31srIZno7X0DnHiTnb04VufjQDuZAZSJvAE
TF9aPiVy+5Cooo0WZSqCs/Qt+AogTDB/lJvkZ2naRzQOO89IpdYQ6dWi5qLd2O5pH4A9SzFJudWO
YbRZ7q+uyeNLYj+lvukZvWIbDyIaST2g9/ZeUv2dZy3rteznVHelZ19hLCGPrG6TdqwzxaQ1FBFd
zqH6uFAHGBVyeyFz7acZz6wEkCjJt3tkF8QqHmmSwOfuEHwvshT2Mw2sJx5WSYI/T36DRDQhbsvx
VTwPkNe+gGLbQtuPMCmW9ym8/2N6xx5yt40H8tXrQOt/noCXx9TJ0WuDJ5j/16ch7g7XUFeRKveB
BNrBnnETnFUmYdN20ojNaOF+2qy/6y6E7sNod3c904FpeZjcr7YJ6imfc9LcMQDHyj3SfuEk+asB
HYEOF88pfiCMEPDOJwn7l8uO1hYPyyfRQtFwMefTgpwNFim+Dbz/RjUfGNr4+ul4e6vCj7gvjYtO
NEuDkj8hvSPRmZA9KFtqb8tX16euIXjATFAosD79LXUnWf/bY0ZvcARgr81I12NVDDRRyvGCnsVu
LQAvDF4SwCW3OmC5MxB0Enox8XNinI5ZrxNglemJo3q8/tipfD6wIwhAsdTBCOcHRIthEgNCcGil
YfgEcAcORQmnxHhCt1xv/oSPKpRnryQ/MlNqTWtW0grDe0TXfbnBiQQdWHg4kyMLAIh0OIAxZrek
nPnrd5ECebPj/PPS8VmFb82b6KuJqDxIQoi3kXRzO2Znf2/XzoLamM5k5d801Kvxvpn8TG1hLCgk
QjEbMx5R4x4XakTnsKWzrGtEe76D79u+e5FXpP3K7Zj3hiF2cZp+DLe8vD08Rl/yt1A2UFa0qRPn
ZpgJ99WLH359QStN2w4Evzc74HEaIjF4BSIHTGcGsYOvYuOroN6og0OeF217SMpdQeaQ5kbT0H4b
5Zdq6MZesBSnVrz3298WkTe7S7GgvGr6+DSPK7yPtRyFS2P0NO0GtAQCgMqvBf1XvKe1LoLXcmyF
UeIIqjghxQ2SwTpDYxGQfc8e8AGGI8JQu7gSDrumDFT0p3nktRyz080EE2W35iQIPTqJmFYg26tW
uQwcnqZu9UHAKeNPkiRuto5gzwYsxkfwov+eT0i/M5cN7aopP5ECnXIK6T+Q/C0K+OrTfqJvmpAk
yl3v03BQL88soL4ks6AEo13AxQQMNCrZPQXaHfX1e2vz7AT32MbQwaApvGQk14+mzhGIfqprz749
llczIoMkpd9zZ+ujIScsjCVI1u9jJEdmAb/PNYVrhyw4aVS1iX56ArvnPoNfqz7mUCSwNc7uO7tv
kZqcyoti4qhsG6QpOD2Zt+pvbpFscpzA0dtpjbSiYvZ2l86C29KjOybCApM86c5CLMnJl5NUdeuf
lZwetV67Fvf+MFOWpa+rCVUmK9oGnX8ZA8iNmigxS5OFbAjNZcZpfLrISl+IjcmfEC2fEv1euuqQ
k3EbiCFkjLi8bb/C9cxZaPH+Hl/ssr/AsU9h+SJJ+H8VnzdotSBZLlVXXVCiCZhAKW0qdDiANKSX
fDmgL4t5pFRIpvoy3yes+JhybvMpuQOJAUL428tUSXZrGX+FQGGmvYo6F5U73Pk4RR48eVxXoLUX
C/SSFgR8dXcTaF3cLsS2zgJuEBexpU3MjuyjhuG3E0jO6Yn8QZmlEC80OQzoNhO1v6acz7iFx4UZ
hkRWqBA8sdrwkOkrLF5Yqlurcu4rvtZANBjP3e5dvEz6JYVHZeuonJMX7t6cfjMXwhq7nfiE2b7N
oly9m8RAXJzxq1h3y6kMA5+jMq0r6JFCDicGtncxWvyosaExvgmIPCCODqbn6FPY5Q3p9sG+d+xh
aumsryXnCOaTr6oCrhEJtmlpUu/K0BhSng9r1XpWFCBgtktCpWALun0kAVkhYPrxgQ3udmVwrBHK
wT7xdQj4FXegDxdfJ/lr28S8IpIsrqwqK0mlKkKzOUQLzALK8PAT5q51NaNoop4ERD5hEIIkp8Br
fKYdLqVjw80HroKU/5h6PtVOrEBuYYQPIAT6Yu8V7oqzCjj9pC5SXpLsHmyh0siKegaGqnEi2KCO
WtPi87tLjNBStGjCSM5aCD/mJr48psp0A7K5YwxAJbb2vyzaDlkLho1tNqMmWboDFlqRP8xKNzqP
d7EIwJgpFtizCB/Zu69sxYMQgOWqR4yD4Ic3vISdON14sSnwtQ0NL2bOEz8z+C65rX6UYxfeM7OY
uxy5AsNflv2cOHo3SVi77vEpEYFrjayRyvu48tjCcVVTKqth+cu64KBLtJcjTMuyD1p0TsTX0hXM
aVKeQrIC5HcPHTgK8i733fBFDOyFcACV9dQ90UaqPVndHhEb5lGaVodzXeiYtn8xUkJxY++upZOy
dABRqJYWGZ8akLMSsJ+73DhvlhSJxlilKkgR4oFa98/VoiN0Tm0F9kWG9SleINlYUakjmz+tuQuJ
a3EcqLzLzf3dAf60+wypk1H9OKSaVJdikYFCwuW/cs5X+KWLE6q93OMvfJVg0i4BCX5T296HajPg
PZLIxYvZLIkF265GOE8F2ASoKN/p019erVl8AbPiJ4gOLRB11qytJCz7G6FmXb41+GgXtGur5xCk
lCZOV0eMabf0Ty3YkeOV/r1yiG7wRjn3Erb7Voaf6u9z24mD/YwWXDL7XpBlTDcVMpLwt9Dn+ZZC
Na8ploc28fzUaTz858BZ1eCEZchguE/f1MOSWbqDItveMwM8SnybBnZ+APksJDKsdRE+z9sL5b+2
vkpnpUJeFoF5SYGa51NO5q3mu/BjzImE0yBR12S6QixzfO+mUOViCEy82O+Hm7YDzgZLu+HkbUgT
a0Y+zcB0JpDQpkOctXwQVslihTB/4UZQTEt5kXkxReusMb6kJi6YgL0tFKzaacbmRSKsamh8beGY
jApXnDuqlYqCMfM3arnTy15qDb/E5z+ON6AaEpU33TAwBWvRFqj1ONFCqaSP2ymRMo0wboTnc3R0
Rg3ZKNWCrTsh1x01VTx7caAbGA95dbd9JFiiTn9kt7U6vStWvttWDuFD7oUgEI6v7T9vU6qvCgHS
XZTFo4vCwcx6zBW+vn5pZOA63VF0jlJnW5jKz2eADUvmTOmqH0vqPvHf8g3/jW1VZBwswGrjJsjc
Q/M9mDjMNcf01LstoR3OwOgaIuSOrQGt1mu/4eHEufyglNZ4hROPBF1USCetLRALY2a5fNypbZpH
nRpG+P8YN4OsFyZEWOcLziVMTFK9qlocJeCyondlQIPodyD+48/EI4wXhUg2wy97ABRhB9IlCGxD
I4xBnEyzRFIhXeWYVojcb2eZuVtWX/tCEiTDaN7LCykqgCWygYoWs/D4kT6uM1JDEFgu+GibdIAz
e+TbYJI4pduNASzLqUjYn4HAVwh54FUMef0fmxMy8aQpCdP9q0nNlSzGuJU9e/gDzNbAb8SeKzDq
c28aicb1TEshEPfdYR0nQ5Sq2XFNbEt5poYHXsk3Fq2uQ5VpHZZVb+lESc64SkTNcJPFpzRaQEaU
o7VnX7QVs4SaSnpaHNmTZozlQxsFsFxZWHZnIaBZ4xNMM4qYgK5ZVnA5cpiK2CDiPIPbhU5MWYKW
PJ5CGbi7nL70Fk19QpZa3kIIwhIkCe7t1y6Lcchkf5VFAlAFzDUWor+hkcySpiU5v69V9Y8ZZoAo
OGqt8FACKOvuIMuLJOkI/xnweiEQQ0Pp/eVyHc5X28/hWs9kYJrT4jXWJiUarDkAz8OMpt7PBBZ/
20spzPkgtm6no4D1E9dioJbPXO5tsjdXxcK6+u33iehj2nJOAZ3G11/Rk0McRMhu/ilalecG6RjE
39cuoI9ji3/lbT++sc6YS/oWJr0iIyZ0R8zGFN05OK038TDxtqpUgKsHEEKWvyt6CX79H+cWGWtc
oSzoQTP26Mqcu6CPxPUlWJCE33916WtpI9WBCzu8niYeuQiqtfepoMud8tolaDmPmic6m1fKA58B
z9pME1aGyWRwpbnoiygp6k/Vm+wPCX86Lfkgzt2cHql0153P27ezpyt/cwuZRU3v39+AVlYMxOnd
oHmsOlcopz5CmiwvKqoVsp1IKaKPWXkveg/kOAw6utXwzL69TyrD+hw6GK4gy1AX6niymS6XTXO7
L1sXsGiJZsPMh2kK/EwjWm8URSx9uLbqJm1Jij+LoibMJpeTARcSPQ+RFzxrXE2D9T7nK8EjGvCT
ecPHxDF8A+zM3jf9U2+JsrXvJy/m2yl1I2f3WZzMow9E9N6VcEJJ3vwc1VxD1yx7LQbN+a/VTUJS
ZK2TrRjil39mseIqJ16fAH0xR5FaeHpa00hgNWOtxv65o+7WHBCUTR4Jsi1vQVpcAo+F2p0QwtE6
U7gUEKNCQT3yDpVn26wiMAJgfXmXMhpWnz2fWQVw91GobYGAW+aXGFcJ1EIt39q/R/tUeS7n66BU
1UDRrhvFBV+JHgVAC6gALXcLJyinA/NY+W0ThD5QHUCmZ2I5vZPtHNztYmc6JBfAJ34+As4XDJs9
OV6qxPhsGfg3vnQ90yToMA1BvVH+qzyxuFuw30byI6byyqt2XrAW1xjW4t5OnHAkz5J0Hb42CQoS
OOq7LqZq0jheSZ/4syJnyDxXrzywEX8VBSLyYVrOUEPcAOAvICCpGs1Vwju9H8PJbE0ctd0jbIvw
e0+M2PY9tuGnU7v5/vbd5aQHca8yljyNj65xywu6qNvPu+VBpgQx7Mc64MEvQHHBhaiOmUkYyA/7
z6gem+0UCTrieqWCl+12TuzMoHH70p4psMoL0iFNCc9LyhpMSi1IbDs8YTrhdrp9yMDvkPaIdH3K
PrBNctdRaLg17q70esMToeATCxH8DJjtQFnjdk1tuoB9a1uAYfu607vBQv+8z0wxGTxEc1aMf7ct
uImMHsKrFxljoouBkQd7GaiSkVsLz/Pozrt5qtrel9pbRKY/Zkwo21i4rSfI9hXzyfrS7ydfZXX1
oHh2y9RFbSSuXtZWjInCqhM3QHfA9Q/Hb9uUdJEfORjHmWKGZu37+Gg3nODx90AiqqkWXDcy8nQB
Ax/hMCqSh0uxyCjLTaYZ7Au37+qa3kqW7QFWQUwbUaYf6PEo6GKEZ18EVzcvh1IuEkT8TWgkwvfB
CD0ZsqhknqCzIMZ6cCxpfYhPtTdaURT4ixyHJLOsa7Bg+x2lgfBxXEwnP/xGbBjm3dWax3RPgwBG
Xa/o1lpt5tXZBGFpSq3coFNqocsOuxRLT1j3RZfEjLHcQ5vWw4y3jMzkiToUaqgPXvbFzhfAu1OI
TER5vPr3v7Jg44FuVP3MnRTmb+8qu6lcP/9cLlQJ4BY37ahKNARwzw+Tsx0InR1uHq0wG6SA2dZ5
jXmqHM5xFYUBKVQf07N8VLw7dtmjqRw0mVUu27IHQsFhTaYNh0pnFoiEyc8Bw6rvn402ihKrn8ES
DAN7NlJX5YeE/mdHqO4IGl3dsC0hvcz65Z78KTazfeDUcYqfgS/BM9d274KPe85fdNmdr1jQC0U4
CY+I8A2upB+/72/r/QYKrZoz0hdinoa0X9/YjSpQ9XEeLZq/t7WFoNAzpphZvSCNUAmng1xSq5oo
ZtQznsP/CRfpcRafbfIPtmQworLMSX+H8+hy3thi40NIFzKeto0/K1oQerOxpueoFeYDEVic99j0
480nAw1klFRtRDeV31/ojzbplpYEEhzYVEDgk/4SUW8ohCMJsRQKOk9JEyIapOUGZwdwpy5UEQQS
uoFXcf1TVrAzwXKeuCPsj92x+jqZsgwRR5A7rKl+aghXJzTir8I8qSZ1swmSurp0wKjkSpaskTH4
EsvZJpIiMIwKkMjdpucwlUw4LwW3Qi/iHrk5KAbM5A/xY/REoqPQx9Ydio0yKjbp6V2sbYzG1A6p
ZMgoz/AArF+9CgjnSRPxVOk+S8oUsq/M7Liy7ry9r54nEiLKf16CHeva01y8Nnqb22GMTe6rHbZQ
ADpttgdS+betw0CJT5CQfHAhnZ3Ez3P0Wg5sVIhtGoEaz+IA30lU/aep1USO12ISLJOcCBOGpzsi
X5tA69UKEWuFjGIMCdnIFpnm+Snsja1g8DR55GANcgDyyYPLnc/lh1SUkOp207KVbkRFYBykeMoQ
WaILW7SUJncG/VUhZ2aCZTMpmNCVKfnQr3B9Cs6y1sJBGzpNqxPJC+23JwqA1ducQaMpH77rO/3b
+5f5s0yrY855LVbatWTkewk5ZlMVC2VvsIvlNeH8RAan1A+ZPOM3kCSBuIezKxNixn9ZS2w2GzE2
/EaMuSvkHWHDAsgi+0e+AOvrgn7Q6aVU+h1QXjE2XlCfb0U60UzUaDfXX+5cKZRygsgKAYGPOZCu
EzWoehLVunPMV2qHp+mjNObu9UV8iwBJ7mGWkQTwiyis0snALGyu/J9C0ybv/yxOjoXx1HHwigAU
FU+NtLz6DKbDI8mKBc2so6jK81CFCoEg9SmAxmUBBVcjJgGUqDw4VXPT8/J4pUDQkbDOB+xGkJhZ
KWR+kofVelQuQgk2PVnBj9kUADejBjAbg6HiXpXjfgkLaQ2sFPB+vyIhILhUN8wpB3VdGTUB4mKG
WnMMoxxkV+JjwKTJI1p6i3uVOnCaXr1wjRGrkVsUjyl2k8ihql0cRIdI/gfMzbwZD2rZJUd3BqLv
DDQlEK2tQwNJpc3FkRPt+THNXbAt44+J+0ZPdjlPTjwq62Sn2G/6WZrLiyPdk93902SptT0EktXw
njCTooNzPj2YqcsAQSHx7L3O+wBfzr+iGRNn7AcWX/nB1YMIy175LW58d57linXDQh1fNdNxCETm
pkhWUPWzQzqPMFnBLx9TEa5FmtjCChNX7Z9jWJy0FUr71JTKvj0IubQVGTbeqrmb2twtStuvBDDm
PuZ3dx2wrOnfcYDh7NpnEJUwQ1Jb6NC22U6s8ZQyYey8l4HeYdsohzmJJLEqijO8WpHtieqjYkz2
UGrbfGMHfqJ2ww7F9ExSgOPuO7XDNYKQQBkYMLfPRKUqYZ1eHpCSDWgfQ5DCRB1HUVqr6Zoq8Qq1
BkAYMPYOerjTii4HuQyRUPZDXoJwWKU3QX8jh/gad7VLQj+6DiUmaXyL+IgJ9xD6fA/cbknZrLHh
ze7NT+0Yhe5jLLxw7IWNSECL2FZlrooGkoY5UHO5u6ziEjdvjev7jZh4ZwB+lhfUJvFjPDm0Z98T
nzGRj3uWvZcCf6GDaRQjMsY6Ptsfz0nZbMHkIvoHCkI0QGpar7fii8wC6/Uzt8E1KxJK/OSlLSzO
0oyeUj/w3rxl5IP2oBNrDtMbuc0ADaPnKVx3XqIJc6Phmjomlchmebrr23nRa0KBtHd9gD7QJy8F
ZXTi+0pOZTBY8Tu4XJkT0Sf2orp4fddzPgQiJcJ/qQhpTZ/CVwveAGW+5ld+8yOfRtRjAtDYfVu0
+86vkj+A2ifH1u6OsvCqgTeB+sItpN7tMrYEHvQqXkAiTQHdlwL4KNAEQCDPzUpg4MqHfDegE87a
KUjzuoWQEzA6AddQ08NTOSmVDadCqoLtu6ifU7U2le2/tLdC5Mx2p6sr/WZXHlJMp5hgvWzbLZiZ
J8xzDV/U1LPigU/LlTxu+KfV6316ZJMNlN3h2mrrtcuomrm3THKN5IfefCa2lfO5JedIE9OMoTg/
YF9PvyoG9B/vJGQRaZ5H/3xiVrVGTxOLQBu0BTz2y6GIAtZN1wdmsfr3IVFqaAEr2i6vAi087OJN
T4+IOLDemuJKmWAXyUAfGcQfz98CoaF9ZAyDU6irRhwKEeS2NCRhi+6tCxbpFCygxKc6xTY/qh6m
C+zhACtzV3fbiy9Eo8t/Su+a/na8nT6K+R3G8k33BkxuWBZQKAp3PVJ8vtOEsUsE2JrcWRzhZp5O
JrTpcPsSUXcF1pb80gQqJtSr5DM+Yw6k1X8+VGy3IhjVXISG81UeAe6UBxLvfEVvHjgcRzZ8CxYK
Ta7ht8PqOPBGoi+osrbFBfkl+ChCyL/zu61z/pQ7zZuOnvST7IEAeg552xGj5zwtmT4lRYkCPvrg
0b+cy/Q5TxntknGaAhI6POW/SssweCLZK6bF1TCGSbrqusp/goTH0QrQFfpRzjRZWUKm8YuYBvvg
CSLNYEfwJyXj16PFxQQnm71zaIysok0cWC2xGasSS1verSy9EqUMG5t3yPAM+niVPsE/VnqkKQ75
7JbKkIB5wPYIvahs8OjSBp+j3jA/heMJSSDjHmDu21Z/4CpnY6ENY6hetyoPVmusD2nIfqzwEnm6
OBKlgITh5j/ImO8zDe286WI0YORY0+C5D0nRcEC7Qw45m8eayJWxtQAukqeSRcf+ejtX8eIoGBPt
brUmlhxKQ1Le78nffPvDpf4BEPFTY/TrNAN57MekqdmIjDPU41R3DU6u5yye0HPxi+/He9AYBD9d
whfIqBieOkL99b2yliFs1r8KegjDjBU3JA7/CRWdH/QyjdO2oOjzHfi2jHoDFgs5DdwQron0Zkgb
BmSqiEhQuzZBNKELcV2TQP+hTqMD/AOHHzOhxUgQ8JMCkzngs9TdPIBYd+zFPudHxiU1R3A886RP
owe7a0aIyEsg9sDnnhBOzD17cZ2lhtwcZA/2SEUs7XIDPGyxnshQSSaRaMJrlFy2SeFBXE0RiX/t
jrsiHtBK4Ni9tIrfrXLMCsA8qVwKd1VrXQthUl0SPYGIOU1dsXO6H6bihDn8rBPDD5UIk93x1njK
i2+9zNsXYqQ9Km7vZ/vnSQ1VoiJUuUoOoXWSGOwKtCsuUoh2g0yHvjClD8E8J6nIzx8UDRA0BST5
zVVGIUFYTnlZ/IaQZZYbpvBqReIzfuyVA1UJAMe3htQlBY/8YPRA+hTEnXgi3NPcZVRnspGHQAZA
Y529uAhqw79C/w8HUOB0btA/UxhtePhqq5xBGdJ4fVQDDEViAWQAsoibseAfgKbRKM3yeS9nm7w4
68N1zaCTMdqRoEUQN0z/PnMXhfIN289+8a/JAMg6Rk7yJbN+/Gw1xdlDiUEIvyMFF4+WFc0MXwxw
XVrfgQGLnll568S8P8cjN6ie9yxrWs+ftocX5X1aa9/QcQX35FhYzXfqdy3ynL+iAwfBGPjAuUPs
SZKFw555K4XAwFd7W2nUeW3nqt1Az+fi3eamBjWT/TNZOXtqbjFWdWVfLufWBQYShNz0BlHbBNQG
5L/3Cuz8imdK/3y1xvywfVAqYFfiUCfq/aSWBH0svL2M0icSbnx46adOT+lbIyaYK5DJ3RENoCZw
XzJmSIEtnCYFOVO2JUSQDo6FcZGRtOjO6ECbF8zFfboFWCerZYu+S/0FlGTKtIoq5nwz3LgKjHrR
7PWvrUUNcQ7DONZp5wghF5Sy6VKyVaEbwDqc75I+yWWyxa4V8wgbkxiLutMiFfdJMUXrTlKEadNR
k2bSeJdH51hvufWeXwrTSL5Vas4wcnTQcQjfHDt8KdIs6dUrg46oQtc3NqB3DiDhBp02BvRLxPf6
r88CcC2eS4OzF4IeTX0+uso4p0ojhM4KqeR5wbaOie3XFF8PTXJGkZNdDSiaPbN2rPn2w8EblWr/
QRyIb178ik1tN+S8xcvsil6jyRbWDFaR0pYX5sKtHRvm27+ClkH8jAyd94Lxs2nHqdiH1ym61LM5
ibaTLawbyrbihhxqUfcGcYyFIpZMCMj6ddHNUIoCCEr/Z9Ly8paHWOUeOzsHD4ofS/d16PQ1nvcN
PMVPM7SOydYDArz9I/OvmRRoqtipmlqayMAaYbMQ2Wi0b/4bvR9K6xjF+R0LGlJIdo6Delg4ehhQ
nDL7GRrr7EsMTwhdHLgSna8tVKd0tGu49d240lDAifBwiTrV/bz6oO3vkPWRKBGBfyldnAuYgjft
/GO09IIPZnHtqiPjEJ7lyO9h2ocm0n89NbDoVatOyDkQ397glgTyLND1tZiKTmCoIBr1jT/K24Cq
1Xx8GOzSiraDy+yGYme3sJm6fw30mZFOrFgrErNQiKQpgqhQVT05AZRrT/kvQj1yYsTYRi8TD1Ub
kriE6wmMMF+i56Jz4LX+Mm+w5RAHyP54GbRJxLsX3S94jERVduSnyEbtq2Z0VMyJ7Qfl9oxZPLyS
i12duNOH7ngI9vtPh4jDLzN2DTuscjpSRppJN4NYNlpj7BTCQ1NOcVUzWExUQJ2ijZxKoDezx00P
aTr+EWNUcBazkOBI4Pfbaer7wG2GXYAjK8C4bxTuMwNFEzOMn188+tEXQtF6KSEfatXNx7gH0xjA
1l10JW66ZnZlt5eZPX0zKTaDgGtTl7UMu47lhz/oOUVHjKdX7KOYLFYOGznskKIBdGtNBRbYTn7t
WxBlAbBYHcKAcMufKQUxSWPaV33Dx/fNZI/56CkE5o1OOsxwsMQp5C9Q1zT2PB2ss10a4hBJhXnD
fYozqoGGVv8NhwUyhTssgvVcckHkiE/Cf9dNzX5vfOoaQ7rKBoZOZx4lR0tVVFVJQMcJbGjG3bte
KeWO4T7bBkjhYrS5v0hI01f5eiejVCB1OnRg2DKYu/1MJArc4P6VVFuTUH+GYqIsyNKb17aoTM1z
ZOEvNy3Bhk84Zt8le41AVhW55bsiI/Tr54vN1KBYo5GnbKcCBgkQURhR85VTsHEyRcAeNVc8+EO/
CFVtvQBL7okO34B+dK/w8KwA8ugNEftVTg4sMT9YkGZzATa+SgNbTDUZ5jYZwHdlmW5JqWeqntAb
KH0YvejdgmvZ2Nea8QODEvZ+1thCMkGpKVVx+HvNX1mP2TEi85aKBQyvVK2n8yOCSAdLc0YL5UOb
gBSgAT+JtReASFye6zAwD8tYGwThLhAhz8I1d9HvZTSUEdoav4PB7XwZVVi1D4cUwm6eWg2JMhMR
zYv+/6FbAO2CZMLbggdh8OHYNKKbt8MrHJoe9vWHxIrGlymfZGCI7TbLRE+8RZp0Z0E3Rfb/xzir
NsNBBGVk6dlB0dEnqg2nur2yPOJN22hLENVC/oM/yS1ve/3vqYI9TjNzRBgIn2GRyw4M6PPY5vJg
S+L+UzQeMShfmaceYMG36xowyCkdc3aG50awGQR+uyxqfKxYmivo8vyHYPoyG6lTL0foaiz6wYNa
4Q/In8q365rWCeHTyy0rWErDXvuwIYlKYfdlRyRR+nslHo9Ma5PuN/ksA+RXKZ8pPLLrdNsmNOLT
If6QCiiXjLWDkC5EJWx8Fx3ZqQBKcn8uUSsCyyYumyxBQd0GzJ5KCPbE6ncEazPY+QQuMyMFobtE
lP+5MHIQ14WY40OZ3p8LcgtmCs/szRxv7KgsrCita6qLO1EtwMEXdDnNblCwcOjlHXBJoH7wkXTU
Je/loH2wtOnYa9OdzQtRsYOnzArHrbrEcJaU2TwB++Fp9NGsIjeeermCjjIIEOn++7aLFzRoNUkw
dgJ4TuW2hFnHcWlbhAZWCTO+wCpkdQ1NgVMSypt4cIf+46viRVl7zvZJHQ0biu8NedK/VMqLIZFx
VNfpyyYKfy4/TrrtFzQgE13CGOfd27W1RPbyfn6BwhM1QXUZggPoWnx8wzG4fw5jdAe5WIOsh5tm
D50QvdIAGWSFTkDiUF8Ic8Xsi9cUCNLk5N6eaY8F9rIsAkEYBQP8p18vSPzE9rnEwLuxujpk3vM8
gwzxCkr6VN7Q+p+nIpM8l291aZ08itK/OPxmmkrXZmCs9KpADNiLg23DlGU1lhMX3da72w245yN8
m7NMnNYs82VPc3zamttLjVNy0u5bmd10Qk+hoDP1sWNHGrPtXSOzpZb0vg75A0eXN41kM4IkrjNg
XGGAXhLYQCyQxHOXmHJAvBosgyoO4/tluOMxiIQO1ZZYYLw/mA4nrKFBicZIGWgcgBvYNnmjD6Sm
WHg6RTtlelny9IEIcoEXD4KJuMejWQ49uMZHevGH/PgcNGfu5bcSH3Redd/F+zuh89JQIgDFR6nP
IMWF//G/HO4JRhkiPyAvrIMLYfQMxpVJDtP0BUDniOgnY1Cf2PYYqbAuVighgap8xtd0CslTWo2t
HaODB5G+vqVX/5ruVTqhleAKKWHr4AJ3/lwkoRmtrXil4mGsnvaaUXG2ctzn3vKF3yFYsTx7SdNw
VMR16Wv5zWnOFwlfqCvLHj0mjapHVY2q01hDHOMLXegxr7TZjLbej1upFWBmywgYD/4r5+VrAPNo
1HqKcJ21rdGtuJgUJZlX5L0sZoDyJWBTI+BO/paRimEBL6yYQc/osQQEw5LmdbcCgIbUl36XqAWC
zgzLgwikKtRAwKwp0XPWdtUlBJfJVLjJlcqO5/RoZdXwRJudfESr2tVlzVJ/vY/ABJ9LXZ7oIAaW
Kq9TIy+GVwjNom+T/IPd8wcjk/Ir+g==
`protect end_protected
