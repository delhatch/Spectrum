��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X���_B�v}�8�x�k.��������A�aɸ�%�ndi���s��NC���zi�8�D��X�i��T�4������LN9*�Ч��t���j���n
����2�q��27��4��/�I ���`Zu��'_M�OJ�,ա�����]�p_��Q�}Ä��"`dmxRUv0I҂��b��wO5�M��־�NG��&V9 ��G�rIg�Qtl8��e���^�^&���6�u$*r����̺��N�= �˜�'~��]���JTbu
�z4|���06�Z�Z"��?��[S!ƿ��z;C�5�9�Ǝ��*�@}�J_�k��ǘq�-2T� c�Rѩ%h%��e�飖
���i��+�o�\:hDղ�z�@߹s�`S�0�+t#�k2"�$��a-?� ��Ɉ�IX�ɺa�����H��׼e���e7�DVJj�a!q'O�wk#o���	�ٻ`�լ�x{8�mޓ=8 uѷ�H�ġ��"M�h{��^���MK�z�Y����a`��WX'���Q/�{�]�^׬��/9���ͩ��*�O�2pѥ�<K�{R��� t���/��9��E��]f%�[A���V$�aa$|��M��MH�ua.p^$��Y�Q� t��n��e�A��d����R|7�c�>4�*+>G~�O�4$���}��Z}�ȑ!��UT7�5傤����s��K��*�ޢN�����F�-g�;�b"���R�_��{o����-��̳�#�|@j^K=u��T��UsQ�e-�@��@��"G�� ��Ko��c��K���B�pXJY0��S�0��1�A�_�_L�g��-<��p��/�G ��/v�
�ceبm�]$~o~��g�#@�|�,���h�5�	�� y��������e<"O��%��#����o�5����5춛v�"��P�#g�,k�� ,���kK�9è���t��YI����#�T,�M�@�,v�HB"@{�����#/o��P�S*��OJv>��߽�Ҹކ����׉�S?�܌~^�C�r�C3H4U��C�,�Y��=�aD#z��?m7$ �f|�M1���Y�W ��yϴ��{�ě�=��{�X��3 �}���K��0�ܴ��TA�O��*��h-���
`̯��Aj��Yn<%��T���4�;�Y��^�@��}7����na5,h�N���o&�_��<ST|��誟?��=]����h֒��vOɗ:ʪKg�4M�0n��nص�c|���:���'A�ь�1(�sĢ3�q'F$8����J�o+k`հ�/Lf��e�kzDe�I���h���IF�ѩ�h��]#<Oa
�g�^��J�qx �0&Z��d;��ڋX�P!;�;����T��m:j��dv���n��Y��˗����������F��Q���q�w�Q�a��A<��o�$�w��Rm�#!+]!�PEy�_<�̏�V�N��Y����Fҭ��pj)�d�t'�L[��t`ӆy�ͩO޻-ct�B��lBa$`�|��)���(��+��Ee#sYkn��Gжu��/����ft���Z,~b��ub��07����)Fl_�;�ެ^����Io�����(�8���a5�����'!�@�6G QfMFh���9�UB#_Y9���B�~��Nr��7��v����P�b�Ҏ������`a�<;կ�tŢ	Η��D9i2����� b��U%�3%N-W�|cAJ�q�|�}۽�~��_j�y���}ޯ@�����$4^�I�j]K���W�����C�vbL��4�|�㷌du���iɏ!�1�?�k�5����5�!m�	q��Cbݺg>���'Mqk9/�yga�v�X"�x1�	���zYz�L��	2�����a��+>X�R���A��*����L/�S:oR��X��$5�<���uWM3=z���O�'~��W���'7Cm��4���p���	����!G,��늁
��R�i�y9�RR���~�
v��������N��֚�Wi<.c������q�X��t�Z��Zd�pO���	 ���Cev@��ecw�E�,��Ӡ�x��5y�7�Wbs4�>W����h�<MrU�1m�^	�����$d5Z��\�b� E~���O���U���ۺ%��C��V�����6�̪���(�mq֧6��9�Z�woF����LK
������J�	�&}e�|���@�DHo��?�d����U�HO9�Q�3�2b�I������s�B5�+ڷ«ae��ؠ���Qp]?�cҷ����T�U�-���#����ӌ�E-�*Lw\���-���5��=_�g)$D<�["ԉ�4j�VB��*��ޟ��B�°�ļ��0��gQK����%����6X�x�Yִj�G)X��[�Qo%�`����һLf������a�iX�\�_�X�QV�n
�e��G�K|t,<�R�V�d(���9&���AN���}�Z���|�{-pwۤ{/�J�V��Ճ�yA�_^&=U�+h�d�Of��f�g�i��xd���}�u>��m���q0�w��~HM �����X��O}�Q['re,�'U��H��E2` sީ�F�?�M�Gj㬺�Z�w�xzs�
Mb?i���-��UB+�]�(A�V�-|�ӄ�,*zz�`�=�en��{Z�6L�c=�4�ïS��yJ^Q�>z�2�	K�z_*AL��a��ej)�O�"��"��Nfr�\3��]W��{�jZ
}��D��Xp�֍:�g��' s��[[�P(�(S#�*��e"� h�\t�U�@U�t��՘v�%- ����-�_�y�nA
�o��&�takiR��c=q���B���٘/��e�!ŲĲ�o�\�nRd̴"��]PO�ʯ�D��K\f������>޽
�PH�I���F��)�9\���wf78]���ģ�ihm!o��o��c�e���0Hc_N.-���	���Q9L%�)�h#��3�q�W�r����:B����?ȶ|�T^zOs�L̩���+�����.��<�Vd&��6Gw�S)��.�M��QL��C� ��X��o��$*Kҙ�m�c�ip��$��Ȇ�����hY��q U{�Ÿ���:i�V�Se�}�~+�����˳�RP�{h ��J8�#b\wu����&��Q�}���zd{g�2Q�x���?��Yf���ꤞt��e$^{��Bs�5��es��T`������������g��J/2�%\�$bER�C���(vt�����>��ûKQD}ι�3�z
���5�ߍ4���H	jI���E0_�-�~0��ۈCb���}h��K�_�!���F.*����Dcy؀)C����i0���
�z�r�������z�<��燱�%����վ"�����R"kĉ��F�b�pch`�9���tLu���k��u�A>�~*"O����}��e4��WB� SI9�k�t�G4���=%���%�Tq�t��#��Q!��9�^*�yB:+�y1���G���C.,�1@��*��3�Y��!䩬�ho��T��e��}o�N0�����$	�����F�*�y2��_G��I쉝�i��=6/
bUF��@�X��˗�P��l�!l�a5Fp4��~�$�nˑ�������9��_����}(g�1]�s��oij!ޠ���C2�N`���`	{ް��t��2o;t���T���qe�1Y/���y�'�&�Oœ��|&�!߶Q�����,���ߕSΞ1�#�I��<����W�g�j~5[tĖ�1|�H�PÐ�s���H��֚��a��d�ݧ"���syy&��A������j'����1O�	�u�M1��n��ӻ�Ɏ,�Y��
�llW�t�
��`{f�`�N�~s�h�-�Z�$�53��|�8$zM( �Z?߈D�����q?��������a���y�7&���r�P�?
c�����+�e�,��?B8B(�c��7�J$i]�����P;�)'����ȩ�vl��I�-�);�����~䮓A�\���e�$�
�N�5~��IӐB�R�I�Z��w򟋠z�j�w�/;S����C9֑�D2�[��?�3����g���h�����`]Qv�-�DΫN�_�ᅽ[_���2r�)�0�n����b�1������A�h3�f�K�ē(������!�9b�n�[FƎ�]��WN\�����fM�W�A�1*_��,.�����]'�}��ދ��,a�Fv�AHj
��;�y�$����Я�e	�f>I�Bhi�۾��)�u"���4d�-Cu�?{��Z:��xܜ)�W�i?#V��k�|A� @�6����	�xT2`�1Lz�7���Y�K�'�]��&̻�.��z�U���Y3
F��FVΔ�.�Zl�ŭN�摬����Y�)P���{��)�㦼!�-h,a���<۱���zL*!E:�N%���N=]{v��ծ���=8�	�~Ov�M�\A$]��6��(�L}(���
��Gk�5����Z��C�:��>��v�a���2�V!�+�u��&y4�*2���q(�C��8�aY�T��ہ^q\�*�So���JO�#���+�m���Fё�o���?-5&o>�I%�6�����!���q�X'9�D2$X?����}�x��;G%(v�ڈ'�p����״?���4�@U%�xPN��`���R�^&q��(��ѽ��~�y��l�1�?���N�*s	�Ɇ�L�������[	�h
�펊��Q9�܆���n.6�Bh���<�Ӯ?��!㢑S0,���VYN�����Z
f:���E6�2p��JG�s���V�g�%����a#��w�|c�t��~���h�6bW��Sr�ya����C���-J�w*΄zJ���վ:O�\�f�+���ܼ���p?A�HyT^�=��OE��L�Pҭ(!F6]Y�@��Z�fv�v�z�*�!��6�69}H�N��PTa�Ť�B�;����N�`���;Cf޽z�L�K�[I����P*����#�@ɛ�7*�.y�|>��mWk8�����D�=m�:\��q$f
���_�;4 �闷����wr|6-��k�0�ku��[�p�W6�Ћ1"����]C	���;`�XQdy��+���JR����ܼ�
e�+���Y�|�[oy$��H���"+W����ʹ	�{�*�FԼ��.�&Ii��)�EZ2��/�Y��9��[��ksb봰�,��Ə�s\�.��ꐄ���tm���`p�����
.%� b�,�z?��N�C�� E+��5Ȅ���ti���,�y��vB>��h��}NO��#lz���#3D�n��B�_[��QuE��{���*��"D&�ÁV0�S��ʵ�D��C�Hs�EtBcpz��4	'��MgqE����oc�U��N���3y�N2w��ô�ܝY���^��$0	����e�/I��5x��`�b(=��B��V,d��i��VY~gCx�}~J��T��q�߀�#��P���x�X~����0�@�3� �!-��$K�z~�f��p�.����m<<c6E��A)����8[�5.c�����o'W��k��Q�t{�XX<�/uZW��0ɺ�J��-c��^o��P���6��ԁɡV����\�ˋ�QU`� y;䅗�珄�B�`�4�1�C߇�xV�e\ķd��� �P�";xR�VPT��5P�Sʛ��i1�SA�6��N��%^�G(�מ;_��aF�]��nV8u��יP�S�6�	Z"R�7��a�vI�m��yx+~��no��97��F×x|:\�"t�?RE]�F��^�鄩F��H�"~��h�| +DW>��]~)�m����6�ծ�󿹕���-Cp�|l�-k�o��^�hQ��ﺍ4-<�}Maz�}k�C����g5�]�;w.�Z(��[:��Y��\SfL�7���E jI��s�I:���J{�!���z��҂�N�$@�O�4�S�p^{�GOCqt�Q#Į${�f}�FՔ���,��\|	T����4ҧ���2r6�Z��!�
nr���٭ͦs̘�����1H��A�Nku��e"��x�s���Ɛo���ʟ�+Kא�=�N�$��j�(0��	i8��ݬ��G W��OLj�������*�[�E����'oWs���O��0�D*��|f�3gT���T�'h��`.T�c��y��0�u��d�5�c.������KK���)8߼Y�%��/~��@&�y(�ٵ�g�쉤�其SW:b����nPC���y���������:����/��^[č�/�J 	���=8�/e���+�շ��TYf�[߆j�+��iv��͐)�m�/m�N!�/,O8w�.o7���f�M�OP²�Vp#���4zZ�5��j0��0Ǣn�B�{���[�{�&��_H�$hU^�s����_Ǖ.�i�A�y6Y*U�����#sW�Ȯ�p�?�]!|��p�u�s�����7\��t^[�uX�Q���V��dO���lq��e�|�x\�Qso���^Ŗ�Σ���[ExU�/�<kQ���F�})F� ��nM���,�%4�Dy�
��z�l�ui�S��#��i��^j��pb���Hm}悚n����tNQ0�z�5�H���Q�$�$����Қg�S�vi����LG��/�|���1���-@2-�A�\g�H���s��K�����)H��C88�����R�D^A�,z�#a�'��X����1S �+�#��6�y'�<�F/Y�#�/�.ݢ���R9(>�T��YbZ�Ui�!��3`&#��r�ۆO-�8QH���W��X��j%"�O�5
6x0"�<��C��@3A�L��Jt����b�D�US�Y�e~�Hq88C������.�#V�B�	p7�N�Q�?���&����}�W��Kl�F�ɒ.W_���d��]E�(
��fIe���vj��(�����^Hl�u~LΥk�>T�aV�.�a�jz,<k����񄇈Ӣdo�i���t�ÅK.��P3xڔ�7K��E���>���A�^<�8����������Z�����a<�3���W�L��E����wg�g*�O�;�+ �4Ws�)�w4�i�� P��O�=G
|�������r#.�	x��N΃�k@�ѽ.$M1p�ι
P��$tYE)3pc��to�Y��Z\�7v�c�(�ad���Y�,���c����W)N7d�Di�.ִ]ʵP�1�$&�nY�J��sޡð��âp��r�i���T(Cк��f}���zc��Q�ީ�㒟�?��Ƅ���2ĥ��$�SG9��dlF&n��#7c�v�Y����AK&9؋^�9��ot��@,�])'�@� ��x>��tQi50&l��:��W.���b_��~�z�[�*���3O��wD��M8�<69+X��%��,�8� /*�#�6]�$U9Zc���a�U�4���T]j/�iΠ�#5��j�%��S�N�Z��0�To��zg�Le�I�o�v�W]�"-�Jk�F��;e#
��ܮ����,0K~M�D�zIp���
 �Y�|���狺�:�x#�m�m�u�$�gp������ؙ��/����P�hgٮ��t��>�`���OD�Ppv����+����):�����RF��BsG�*�b��W�C5R�u�^�I}�<��C�~��&v��/�YR�ٝ�k.��k1�d��,(G�P��Xm��m�M�S�4��h�xu�'��')M�*!����! ���˚©��w��Lɤ]�;V�~��D�*���|v��	tC�?矀'm���9w������#'1�Ѹ�Hڙ�&�0�=D�~Xk��"o2ح*h�~_l��'�x�<��T�y�3]��͕^mb�p�,�P$i3v���l d����l�l�NF����
��ݻ���`�r;��%t�����kZ�H~X��c��e7�L��n�����[�T��y}��K5�;a�����#��+v�I��q�3�����3��z�]?��X�?f���!��~�d�A�we=sސ��j�K�<%�a�E��=�mv��oj(f�p��=G�@�� c����̦t��[���4�������7�p�it�Զ�����{�i�p�B��;�~-�V�G�!�� �#����8ݟH\��Y�l��-���*�{=��궙x����6��W��u��Ù'O�L�����2h��rl����~N�f���$��<ܺ<�tcX�ݗa����K�lR*�8�"D@��WTE�M-Ģ���(�ޤ��tq���Y�b���l#j��_��/�7��'.z�P�hJ��i��1��f_zc�`a��(x�|���r�ۗG�����fB�mz/V�E7[�y��HS���@l%��݆�{�ќ`�co_
��v*�uY%�Ψ��kjpV��}�.ǪT���^r��u�ܨ��M��t��H'��WU��%�U�9g{'!�n$8jr4g���=����]�|��L"���Q�ļ�q��_���3#�߅�8Lv|u��@���a���9�fa���,j�fW�n�Ɠ��*�^[i����ny��K.�Bsz=W��x�ZD
�h��O��2�ٛ�1Z���.D�-�kXakg��W���gZm���#T�bힳ��=��
r�)<�ڝ����@��y��u^ؓ�mT�
ܠ�+J<N�"I���
d`L������cNN�S���M�j�j��<s�n�x;4�fD�W�_�������}������Dz��P���F��#e�վ)[!�$S,���ce�?��GR�Q��^��W�F�����2*����#[�p�q�kWK��ƀ�M��^�׆٫���
��,
H�W�R�,�^���;�%����*�x&�-0!�4{ju��`�i�Tm�<��dcwG�li��\��������~���8�����_˫B!�ڞ��O��`��n�����E��V��}ˈ!��z ܝ���
"�ne(J�k��Q���9��$[ﲆv'�H�X���"�-��*�9E���7l	��n�e�J����� Y):k ����+��Qk�}�������of�J����Z5�7nZTs�m}�U��!�~� �߮�3n�l�;���.eQ��5�gF�� ��}u�D
1��5��x�zm40{���}��Y�
P�D������Qb{���X�h�0l[+�B���>CF����jZR������Q�V��r�D��c�_R��[�)��������(y�h*D1�c����$U�=	0#�P��ɟ�n�hş���Y1�A/8h|{�&�T����1��8��Y&%�X�	�5<���JD�eo���BDY��̛��[)�_*��(H[y~e��!Yю�77
�����ß�fu�Fa��͊� �^g�eQ��yJ�����\�GgbK�>ޡ-' 9+b.�]7�x�P�(r��)�j�[�S�p%#M�ľ��CC5^N�B"�6��NK3۞S�}~KSk��2��"�P���--�#"�+�u��|j@x�4��i��〘*��ܭ�NN�j�W*�z����$��^����B����M\�ow�y@��j���aEr]NctT&G�l��*vF��H6��-�7o׫���}&{A��P2���aX�C@��k(�2�{�\�����R�f��'5��-��#���+�R���hĒ�`6�ʬ\���˟��Y`��
��m>g��HKsd����n��3�A�=V�/�q��"�ӄ#@��ʷ��}�	`u�8=I
KG$�����Ȭ�R��U��12�qW-߼_)��vk���`
�Vy[��^���PB7�r��;��0���,`Ѯ��sf��G��{��=��I�02E�?�pR�c'<=��r�#Ҵ�i��&VJ.
�C���+�n_Y�k�W���a$!�-��Ф� �H��L�^��ʫ�T�/���Z>��[/�Y��M�!>�*2_���[":6o}������u��U8��&��m�aK��qBhn^�mͱ�T�N�����������N0�	�O���.	�/.�����Ut�K��U����X��ӳɥ�Kw�|E�4z�u)�\�`�= 'k�x_aL�z�.���:S>�L��	Qa�7Y�U�G.�x�a����;�:>*��sTaE0)/���^����$�h��zq��J-�!������UjmN�By�SaD�;�h)��5��L���TT��OcHGV�rG�Տ�pL�!�va����g��k2�����L����1�>���	t�98���m��pj���
��>d���ns�,�+����Z�X=���7�U�l�"';"��ы!����j&���ͦ�.��`
'8���\!����l�2���F�1�W�G�n����~aY�c�9Q�=�T{��6�{�d^�^�w2+i/+ߡ� ����M���}�T#����k)��o�S_h:e�f�<�`O��	V��Ɠ2&'� �	:?���Z��WK��]���)Qe%"0sј�
Ol<|�H�ᅩފKE���[U-b�w%K9z����(}h,4/e3���Nǣ,Gci�J�?���F�b�hrCrGf'�CvP�v3O�X��Uҩ,�p��q�9���e�B4h�\�t��
��'�b���iM����f5� ���a<���
A󫣄�
�{n��E�3�.UT,Tjh�b։ \���ö-!�Ƭ�#�Vn�WPaMU�!��Ng)���-+R'��T�g6�](&�$a�0�f�t)̃H9���?J�n�O��4'F�E���t�����-q�3�	�8E\��B�	Z���I�gv�^��Rop��Q����'B���7@�����{F���㛖�������� u��O$���$-sK=����vH��z�fq��CV}�Ǐ��y���(:�����,~�/�.-.ce�6�=�/5v�iIg��<⩨3�nv��7�]%�v�Q�a���_ݣ t�$��h����bŎ_��.��Ej��O_ݗ�����a\��X�]�c�JE"OG�ZWP�G�2�{�����&��`�N��vw�Y��"h���6�
�ċ���e���A�.	3;R�E*�Q%�T��e��� K�kw�k>�t�����	�Y�$j�8���c��B�1�����M���4q��o��\�N�0��+
�#�w�YZ�,��ٜL1,����>�\����N��&}ЍZ���V�$��ȗ��}���ɝ�Hel6�V�}W�#c��^Z� !����f]���+��248W�	�͖��_����W�`7���?g�;�-��{	ܖzd!őT7 O���09�iŋp2�� �3���E����A��e�TP�q�\��^^���Ł������"�-	-$��Q��i Y	1���vT�z�`��X`�@Vd�ҳ��~�g���2ګ���DO����,��"��v���:����됆'��#���NH��+}"^�UQ�����u���`%���8[��kɬ�b3%���2]}m�ĺS��7�>ZL�����M@3oJ���<}	���L�9�Q�q;f9n�ύ�*���s��KL^�(>K�z�l��Q)Zefo��崻}%9�)��`�+�Rv�*{�� |�Li��7pҹѴ�������O�-��7P�F�،��U�s��nџ\|��kEAo�
�/����D��tTa���%E�/�C�,oR>��"�G�7��O��;���wY�O'El�v�������>�L������3�k{}��;��y�����e>��tZ&x4Y:}Bl���я\��/� ��T1��( ��LN�
��vA�tA������(�N��=Ph�����B�\0	�k7�f$�ȵ���?�U���`m�sm�V�n`���M�[�'u��=U�\�1j��fj���̦3q��-�!,֎M �}�Y�yr���x � ���;����GDD'}-9�^����֌�sL�U����b)�]�ڟ��YV�oɽ��z���U
��U"�i�'����`z�����M	ON�+��ᵕ�h��t<��ˍ.Z��g��]�{�8날��~����~�0�W�GLr���H�� �֦2
-澞��]����z��R��iM�����LI��n�"Gnק�Z�5�I�`r%�n�$�uuwAդ`�c���o� ���{c���];ϡQ��sY�?��qR��X(��54|���կʾ4ɋ��Ո�,��ۓH{-���җ1���l	3cbϰ9튢�R����\\Ֆa��W��苜�[F1��?Ͱ�7�.���G'�O��H����6{����&+��_�G��Po�>%���g��ڤ�H�5Sd����-�F�]���c 8�����I��xA�K�;Z?�X��9������'�"�vFn;�H�;�(H7����'�W��d��)2�/�굧ο��+BT0/	��>#]���a��1?"���ǉ��8YA���,%��!����*�~Lտ�� %>��2C��IV��W�V[�1�9�1P�Ӏ���2K���Wԩˮ��(,'s��CƮڙ} ���0�8�V7j �){�C�Р4����.�R����_I�[��O��,����,�;IJÌ�a��u� �ѹ�g���rJ��(��@���G����>z:��:���ή�K�$�r�ֹi�]~����=���g;��/��R��Oz���Ծ�
�U�
�y�V��#hL��1M�}��	z<�����޲!e��P>N!�V��+�Yf��3�ج�w��'�㧷7Ż���+t�A1�2F�b�~}H����o��c�]`� �q�*�z�a�\�_���J��ԅ֐>dv���d����ē�(4L�)�6e,��H�D�:�q[:`�q7_Į$١�z@��#,�@�����uf(S��B
�	�\j�љ�WT���[����%W��m�$r&M���H=����]�܋�L~<�ڒ�9��[�tS�k����U\��S�w�1������m�đ}9�UR*!��Eͥ�2E�����Z}��+?{��$l�wo���Tj
��1(k.˸	���).PPr���]B��v��2Y��	i��!JK���
7��������U3�4��(H��n�e�MN��w���"���(X��1�⍑؄v�Ȼ�܁E=���3��N��Ϲ�?�����GE�G�u��o����ohw��-�`�e)�Tn�wH�+�Џ	�F��-�3[[����`�yPl.�L՟�S�Ż	.p��j
�e�s��)Ç���2v}�xDp��#8m`c_��r�DT�>��y`��Q7�V�~m�� �T=�l�����2�Tq|$S�&��)��vW�gg�S�P�>b�ˮT_����J�����j�)�a]ʅڴӓ�
�I�H9C>�'�;9+sT��^ks��CV�|K+�FB5L�D�琟�&%�3y�)?�mv�ҝ��`��ց�Y����6QE��mV����Y<��_�P��s[��b6���ucM���;�`=���}���F�=�y]T�żz!<��<ld0�b��g�J�r�U@#�W�g`�����]re����zf���M�ʺ��?�A�;dq�[W�A��ALb�G�h5L� ��=�{�@�Өx��v��@��<�(�ൊhw h��n�c�%�{��Jx�?_���V|�5��t'�����a��3R�T���]5�@�\��}�089����
�L��l��������/\�/t#̏ ���]�&ML8�_w��$a���m��֎��&8��A% l	3�[a`4� �|��~v�˨�� ����$�EsPH�}�����1CEv|F ��5Q��"�ag0�b2��#p��4���������ޖ8��_�S�,���a}�>e%h���ӭ"A[ ���B�X9�hJ�Fk<ԛ�|?LVYՁB��u���W������������u������x��0.\���>��p�yY(}#wLTۊ�bAkU>��T�MTx�g>�5���E�ǅ򅗘�Q|��%��r�u�Y,C�0�/��_C�o����+7��j��M^cH�� 0���ْ˼�;1���t5��z�L`���?f%�z��8 ���/~^Ŷ>/�?{�&��)b�|���o\č:,���Q�hM�+B`F���݆�Rw�W��HB����d�hC��uk�=�p��A�����+)"��uU�?��ʆPA���+���.�-'�hG��.�b,�CH����4��*GY��?{���&���3b�4�?T�̝�=n"������p�L`fdE�E��;L���9�6&���kDж�ت��|���,`�Vqw�-⻚�_��Z�<pOA���ғ�����8���B.�#u���t����ͭO��)�Wh�qi�pq�]@�a�gN8�q�OT&����t_�	R ���'���Ђ��o%����WnK
~L��?�`���P�f��g8������|��?����޺~�34�>���K��n����㢏�����%�ԭ������%q�m�s-����-���nXY0`�ci���X�5P?\Q��4³j5Tb�w� �s-#e��W�'R|��+-��~�/#"1���)l]@ ���4��c�m�F�|�? f�9�!���o`�0�����E)%
R�	������mv<8��7���'��d���j^�<�!�Ql����V�b��v���3n�, ,T|�����!�|n���M����j�Z'o�@�mc�ŗ`��6Gႚc^��'�v��'�
�j�,�ŉ0"��!��b�:��o�1C�X�sLPB�3-K���ݛ$�%qE���+<�9U�e%R���H"�e�V{H�U�lo1I6z�XÂ0n�۰�e�yȶ�[��G���t]�b�]]5s��QN
u��'lwL]�ztX�s4�ɣZ�DbbN�t�u��#�'%c�:����)�D�0���ǥ{�wb6]_(57�:$��'k�̿���xA��x�xv���Q����*� ���\'뵝�)!>5������as��hv��o -Zw]�#m�YrM�s,�96v�㠵�7�ErP��|a�
���h^�o	��w!��%��I������jz.ӣv�D��Q���H��7d{��[N�����UJ2�B۞�@i�b�I9�t|�)ù�Tr��!�y�V5�ȵ�d��9���i+�͸�P@|5�b����=�_�%!HP�{�Lo���������{��nK�5�x�R�%\*@�)I���l���Jﬠ����m���!�!Ӊ���N����G/����2�R'ް�_��1sC��W,��J���
8C��aZ��[s˽P<�?$6���d�j�΀�|�ąՋRS  ��E�dƋ���yZ�o������dq���ZN]����]�@���P�ن�E���ة�����J� ����]��.�ݶ7�Km�"
=>S�p�+{���s�@)n�K�˼�x�hTd`Ry:\%Ck�۾�+-k"������t�y"0k��BK�\@G�%�&�&OhG.`Mt`�;����o. �1�U�T�S�.?�aF�j�T�Uy�A1����m�G�$�ʣ[ǚ�CE[�����t]�fk���dJH;nz���'���	��Mh�o�7[�'��q��D-�1X�=���J��U����$������c-�������D�^�D2��!��<AgCE��� �����	f;?~z�:��
UH�"d|,n�$1'�z}���'l�\Z/m�#;H���U3�`c+px�i*<.Ԓq�o�Ib�X�_�Ca�l��s��:;9�H}1�=;����
F�f�� ݬ��S[[+���� �}^�%���%s�O�;g
��d�\@�Z�Ҟ�yuX�p��G9T���5�f1��e�s8��٨�}4����=�I��D{ܘ���f�u!��Gm2��A�>�7mrE�M��w{�8���ՙ&��_">\�ֳ�|K3Dғ+7���O�C�A�~}+9@8�9��ǹYQ��v>���{�a7�3����#E*}�k�Oi���c�ݖ؀����8F�`V����r�cA1�@ڌ��S��r�����������z��!^��{&�͡ :?Ov�ːP��m��p����y�~�s�E)�.u`D�q<ϻn6'��n�B�L�X���4�ռC8�,�����5�~�Ȟ/�ʘ�>j���j�N7��1Ǫ����E��QJ]Ǣ�ݸ�@��r��Sh���G�2�Uzz�1�'"�ö��q�0��kZ�D���E���\��}�&��L��=��6�Okط���m��C�{+�@�����r�:3= n��'�2觃N7��s���L��_�Q͓:�b9ݫE����H�MQ�%8*�p���ܔ)k 	l2�.���p벛�J�^	+�,��s���r5���rz<�M�ι��Ԫ�X����]�7����7lMv���>]�E�'� 0���̝���=*:O5��֙��G�^I��x����@R6ڼ)i�������vi�ӟ �/̊�,��i<��Q�*�9��k�z�����S�G��TѴt�0�s����M�kn�#�z����83��a��=���B�)H���:�E��]h�լ��P��K{	-Y���ܽ�@5\�E�+�ȕ��*�3FF�Z�/�e9o�뾋\VGā�ZG�D=���<�5��b��)ѹ��C���mc��x�c�4Z�m]N0�]�G��@57�o�.�=3�c��>{G|Q�lĂ��D��vC�b�皨�
�.���a���6���D�!n��)��p���c�f��e�'3���IXаt;����@��`�R�^E^
ޭAc!gb�x�ع$>��n�?ً��_��&U���$��x
(��c�^#���n�u*oȿ5_�"d��|z�8]V/�� ;�X�������j�j�VN�hg�~l~�Fj��'�Ԋ`����B􏗥�+�牕W��H�s�I���3*:�.����@ N���^UH���`.�a�A6۳g�]@[�4�T&T��z�k�dS��1
�w>����S���*���3ѣF�O�a�W�]�CT#�S8��T.�֡�N0
�)t�ze�f�=^��������/�X�@�KK����U�w{:/!#�Ǣ�PC:/�:�*]�!P�*yn姅�J	�t���2]��I'kU���Оjc���+�tXځ">��߯�r����B_�`
�פ=ځ��"�U�2��R�������*Me�.��h���g�Dߙ�o�-�~��T��f��J��&y}�1QS��z�;���������'6@(� ��`���A�w	3)C�HJ�*�������|�0�Esft�+�M��+Ei���$:40�{�RJZ-�7^�d�$42�DϿ�<_�EX ���aT�LTF
b���B\���^�\)~|@D4�c��$��1`�N*������aV%����G厑�Y0}�N\��,��"��<3xbY�$��S�xi��ݏ����˛�$y�IIب	Y�#mE��N$?�e�o��=m6��u �����{�0&�]��"h��`~�KmPP,��=^�AR�5`��������b3&�6߶DM8b�aṓy��<L��@���ȱ�j?�m]�,R���3��6���W�@��QT�<�\���t	��Z����G��}�HxfjAp��mp�`6A�9M�4����j?Y7��|�*�Ѡ��}If*�T���<���>k��� .�@ޚiD�hq����C�. �\Tݴ�C÷������]q�����!o/~��k�����L�Ӳ�m���0�r�g�j����i�H»9�|h�"Өi?�Hݗ�o걆��tP�I8�Wn��W �y��3��5_DfjF+Y� �������/
P��Y�j�$�׷���R-�����^
]�t��e��u��H-U���k���8<'�g�T[�(|5ޝQ(dEE�KEom]�ł��m��KcS�d��+���
�s%���o+�CŇ �JC�܎_����-��5��V%A��A��x7�2PN��.�o�_�s�NͭN�p�|:�AV14�p�V�����5���ҝy�� ¥�|� ���A����}�'��B�#��;�U��o���x�mxA=e�Ep�� (��fA��B"�S��CФ��R�@���0�7(�ÃTQaMLeוc��oqZ�M�E̴�Q^`a;�W�:��כN�L��n���2���v\��qN@'�g�������|�e��۝��|w8�"��ZZ�bnF{bɭ�6sy�����t�}䐑���~���/�P5p�*�<)%�D�@�)[��"�ݗ�{a@):Ї�v0���!���*r|��ۓzr(�� /�B�0"�uקG�e��pu�o��L���/r�$w��oY�rB���,�
��z�a(����i+ �4�~C�e�Q����z:z��Ə+l�(ZL�6�U�V:�f	&�hqJ�a�毟�h��j{���CNN���u�[��G�F�'�AԞ����H3\�].8&�Z��A��\�z�l,kd��4�3z��Bn�	�N��T����*��r��\N�H�I�Ù�S$e�+Q�6)թ0lO{SIhO;�g�q�w�i��Ya!JJ����OM�+����6���>��aq����O�a&��Ҽ'�b!�xzr Z@��sFU���B���X�1pP<�ul�D(<�e Z�VXG�˻�a��޳�r���:�Z���':�A��
�_uv�f��q��s�Δ ]ei�	6A�陡�G��C�����	���'��L��'$�?��=2,缃�e��J%��E�j���k��%q��IE�/�G���6h���YL���1 �Q�T��!��0��� �2�Wk�<�'-�l��g�A����T'����>�E�g�vv��P�(�h��\SW�t8��� "��l�����G��xU#?�Q�P�/�! M�h������������F/8^����9O ��8T�}������]�F�{�ƈ���'g�u�9��\MD8��V�Z5���2�rJ���6���8�%�M�	�
cPj�A��΂^��s?��:3c�)��3��βJ<1 �sv�z׉�[��ͮW�l�5���5���QH[jX'�k����ҸU��9�}1���L�g��W��_�Ji��C��B�.��$���\�lC��~@��NZ>x��Vé#�Wi�p5,�(~
9��dNP wu���h\��b����hX�'y���;HX���L8�M�	��� ��q�"���~��ƥ����ˮ�Q���� ��uI�K�5x�F���=�:��Y{;�Z�!;Z�� כ�n��(;��h
�h{�Ю��)�2��:y��х��拞�p����������%��0ڕ�2S�3�J_�F� ��{h��Г>C.�J<��<?(c������
�<-�!r�bf��S��- h׷#k��Әu�����^�'\+#�M.n�����d����Я���a�+��/���A��3>cQH'
ܩ�4�	���jڲ�H.׫�����Z� D#���a�ͮ����i�H�@�c�)^�AG�c��b�	X[�BA�o�B���VL��e�y�?�x�E�y_~�~�|�z�p�:�j��ͳ�v|��-JX�Q$u`�;-k'��iYqd��p
�\˹o)?2���F�g�IL_Y��i��#�iЭ�5��Ó��]�GͬK�%��-7�rfzxR$��0���Ur�*Kd�=�WY3�MT���2oH�]Ӛ�!*��TQ�9�Y���Y��z�c]���G2pm�G�xZ�2/���y��GĮ�۝ڔ��H����}+�]v�xR0�y� ���:]^F�_�R�g��ٞ�2�vM:�&�>�` j>�~.�xbZQ6�w��A�V|*��oL^i��n�=Ў�ifX-�Es��B#`,kâ�3���3t9<��³�C�<���1�f&�. �5{��Ʀ���Ύ�cqA��w��w�7��H�X4Z��h��������7po�C�OUd]�m���8)Y���<�LW�j���
c���A`|>�U���x�Zb��А���Q�a��_��J����0�Y��#��.D��z�#M4*�Y$V�@_p�Y��*"LL��C�=�������I>A���;�.`���8o�ۡv�x� '�	t�+��	�.0/�S��º�O����a���s23D�A��H�!Yw�	 �gP,>���"�m��5_��s����\�1���x�8i��d���“���`�H��˽���kU�d�i�^��O�^ O�*v�I�J�wlW��ˁZ����?���^�40�%��ȧ��վ"�'��6!��q9�B��Te]Y���`��T�Z���vX)Z��K�mV?�-4B&��E�x�̨�P�R�V���C���^�c'���	�x*�F�Mł��Ք��'B�H�ۘ_T&��?5@�F���hE�og�.�Y`4��p2E.6���}����%��-*j�ȋ��p
��:��)U� "8�Yw�- Ea:�%��ԇ�#�C�n��~�Uyĩg��cHNp���������V�t��]���q��r�����q�b
��S<>s�[no��Br�p���i�y������Zo��h��-�K�c"�<e.��Fֿ�ߖ���+!�zt"�k#Z���פY�:��v	{@��uJ��ϼD]�qʹ &G Zb$2�� ��#�AdY�{���r޽Z#�<����Ah��>QY @#��4�Xy�n�R@5_%����`��,��jl��5k�b�pY��Z��3��nF�:"Eo{�AVǡ���f�)Ӯyk�i�
��<��H.�g!���	�%;s
��#%�D.1���4�}�\�IN�(�R=��Z��[_��ӆw�;�#*Qv���Z>~�o��4��%�P��}�<�����Eߐށ&��`l������ uq��!̈́�p=Էs{�ָq	���؂�$���~cz�ඡ�	����}ӵ�H-�o�C�ՙ����s����"V�4떱8���"������!�O�*E9$v�W�w�'�@�an�p�>Њ��7�����V}aԖm�#oǘ�h"=J��'C���Q+�3O��{�i�襵�A� ��J����IA���~î�W	u�p��h-�� �N����8pIH%�;�<��۳��8������I�_�g� ������m��yc�4��L�T!pM�`Gz�f�U����j���OP���zQ{.��.�W���A�έ��pP��$�o-���;��f�F.�ps�Q�G8O>��_���l}~0��� 9��@h����KI����̬0���&�xX
�ЦF��z�[������� �j�~��9���o��0�H&p�Ț�(UEjɱ'IY:��>�D>�#ՋOGu�� K���\�F�؞����-l�i��%�����Y�ŕ��)_�=��\ږ��N���U��̫�kS������&�i��k���8��uJˢ�&ٺ�S��P9�s7������F�lW}�.&����?��O�1<Y�"�rb1J�����-��dJ����/\@>�-%�J���dw"��ZZ�P����b⊉کJ���">���L�`_='�r�v�,�Ǖ��%KAn̂p�z'���:-ކ9����|w�T�Ś��)���o�m�^�+�G�=<�OrV	�+Ƀ �B~��
��N�i��i�n)o�.ŕh]Zd+�q3�{{}//#2;������ׇ[�ymNXJDőI�&��
	g��̫C��m�Kn��W�x'���u�qt��)3�mIp�}�9+P�<v6щ7��N.Q�Mb)��v>9�bAm�x7���Ѭ�wd�˸-݊/��\&�B�c�>�,u%-��IvGy@nM��H.N]��,2߈K��i`�����k/-����"��,�p(�Jv��:�btT����f��SA ��^�Df#��|��s߭����;j���S�$>z�ʆ�s�{����.����m���u�m�n$M��/�ӛ���X~�!zۖ�>����^Ҁ��J\&�;d���Ͽ�I�;��Y)��?�0lAM�wn#��'�U��u9#tm)�f_��+[~�s̢����)�w(]\L{d��G���#�TD�\FÒKq�EԪE�[d ���<�4�n�ݩ�p���S١Z����W[CE�y�7D��U!�W��v�H�Qx"�����cI\6�S	&9uRH����f�X<�ڬ�i�b� �b.�Tb�k|�S��\ �a�?������yԹt�8��4�۹��3�k��])¢�j� ��ί�����Tc���(LD�) 
=�׭N�D���J��l������1-�|����qC�+����f��Ѵ}	�C �gy׉YݴW�A�x�4�6]�����"URy��Dٿ�)����1}�-�]��9}1�}Y��Lcn�=t�r̛�V(�x�P��c�� ����KV�&R*�I�\�0d>K��!C��ѱ2��Y˪:^�=+��S#CD��ݙ�x��#f�סՓ�U�p�a�k�|��+FPV�#�O��n!O�~��Q��{Ek�?�D���.q	ff��P�_�O��^��Fk;��*���[�Į�쵼z�5���٣
s�:/`����4PD��>!���5�
���*��I(��{�Y�o#>(S�������j
<͐�hc��R���G&��t�k��d����Qm���f�_Ɯ2b��lhP�M��|� ?����^�|�����넋�vhT8ӗV��q4�-R�-]+�GxΩ�Ttp����x8Zd�a�����`a�{��%�/X�L-���5oHW��Q��*�Q��sрʐE�XO����A����*M���&�N�5��I)���5X]Z~�TC{&����O�0IY��1��Kw����;v+\�;{��o�hf�hȞ��D黆� ���G0:Y�S�B�-��0����m�&��1#�.V;QЅ�8)��5���7�\��	DD�2ɲ��ha��K��z��0=���~RrD�-�w�3�%�TΠ�o Yi�Mޚ��&����o`ۛ��4�c�Y��ằz����8
*/��;>�h'�^���-z���b��2�`�r�E��ӫ� \��>x�U����B{Ɇ�>֨���A� ��GQ��T�O_1-i=cB,��M���Ȯ`��צ ,��� x^�Ćw�w麥j�w� �+m��Y�Uc����6ڟ�F{(�1���2��\5�=y4�8{�ו=�"�R�c��]��V~�h�-�+��4c,�=n�\��Z+��a�È���I��z�)���1��M�	�B���n$��J�^<��J�IX�{�z�֞����D�r�K� (Q@������
��#����;c4�G�{[���E��V>ht wR<9'���#1���ވ��X�qů�Z��%�T)��4H����J�@K��с�2�_&*��&���������o���80���*�f�O㷚��(�`�	eT��V��f�'^�$�o%�AurP��G߂eE_Q	���␋���'��#%��*	��!�� H x[#V�W}��$
h�k��n�H�1C�zp!�A
���,���:���o߼�wcb�5o��z9��c��2E����ᵱxW��E��d�������`�M7�w��U��}H��B@����)�x;<L]�E�Cl�4MjÞ;	���cx^4��9@��˷�~CO`:��/����ly�o���&t�;�����g[�H���6v�BO�ŝ%	�`��;D��6���g�lV���C�B� �N��"<S��Q67$K6��������eswT��=d����'��Za�7B��7��@ݞ^��ͷ��
�&�"�����6m�d��_/"��x��Jr��f�ڰ����D���|Ψ���n��Bi���L�>8eo�A	�G�afO����q��^L�:�Q�3���5����73����y�����%�Q���H��q ��.��X�#�b`o3��
�ԚT1�4~"P��y�̭�+�'UҼ���o�}�e��W�V������*�k�[��t:}��X�IEo��.���R�8��gB��t��B����tk�\� ���	�)�� � vt�p��~�?�2*6?�Y�,��=p^/��{�M����z����̮r�����r
�@��5�p���o���ya���[;���RfHM8���WV���_�=ۘn��Z*b�Տ�Oy:��Na�m@��'�j�P�2����26V4�+\��ܸ̇�/&(���Lo= �ИF>�Ӽt��v>Nt�!�UHuR$eq�b�r-�+���k��At%�=JJ�� ��������9���޳��&W�#�<��m~k�j�͎Q��[�=��k_�Xz�׭��uG̭9\����a#X%=��<j��۞yu�g�"���o�'���b4���)p}X�{ Y�{g[R��3E��]�s���aK*������4v�#��;߬��l�9���6*��x�o��g�S��77��"���~�(�z,���A�@[w�-��D5O�Z��5����u��u��R�tÎ RgH�X���,�"\k��hw7e���R��`����xY��Ěcڨ�,���۾ý�͓�xp��l!k{+�c�;l�����lM7��]��.&�|��M\�x.�������*
��w`��+���[v�֤����Bo�C~l31՝�	Y��M�d'�����(Z��`^ܹ�3s:fѩ���D�=�I�	�K&+a�\C�1�ea����F������L4WD��z~90,Z(F���c(;rZc���;�)PĲ��pR=*��.���.6 r��\I�U��:J�c��6�$��4��\Vk#�o���6�}DG"W��r-N[���SF�e��/ �l��B �}z5��&n�6psK��gQ�D��`�!����Z7;W��f؊���R�0m�F�gT����ᜟʅiSA��1���@����ݚ_|&���H���øQ��f.�\㧖ħjd�)%��T�ɐ^�x�j��C���.꨾oE�p����x�~��@��QZ�k�-��N!( fv
��Q��^dږ	��N��(B�a�aF[��O�
( 
bS�ٚ���5\Jh�?���6�ƈ�BH��{G��oG�*���1��oC��nΤ,�u������ݟh^�
ں�BBAIpT���=�n!f���������&�d�b��1��u�iӽl�u����A���w)	/���
��z��,cw�����_� B��n&��4�S��Z�H��("8�5���EV�co���yꓱ�"���������\�#ڊ�p�����Tq��l@��˳Ƴ���
� n̎(a�9�� �L�R�*����1=S�D��1�e�ڮ�2�銗�z#�G-���@LO��'Wg��UPߓ�`F��@kz5b�;���k%wu�ǃ1�9��39a��lA�H��n�u��*����}���}o1�1x�X�,q~y��Z����]C�+��Zp�a|���Q��5C����R�Gx��
?��9'x��J���lÈ�3�V�6i�Ti�d������u+�.d:O�O#�B���.�h2}ō�2W�=���=	t���~|+�T��ݸ߽0�B�ծKF[�^X�@�6>��������v��1"�J0��X����/��d�:处%�3g�ypXDL�=�ZA�]�#�:m�;|��[��k�%�ߊ�NZ�]�-qqq�S�㩹%��9�_��"�"6�d��+��*σ:��'�~F�˳h'��[ Z!ʦ׉�d)LA�$^;�����~W�dC݉h��Џ��m��晑����^�)R��r�U��c��gKt1�]����T�O��+�!��&�\n?]�nz2]e��nT��v�f�^�%7@/�:���u0J���х�m�W(IGm׶ ��W�pw�#�����;8뮊`���c��Z�nO5"�(TR��,P�%���P6)7�f����`[�y��U�Ҧ�\ �����m�F���[C��?<�췌�2/�_"�*3��5��h�f�-��t�B�E�xK�f.Q���I��bi�񬘱�"�yZԤ�:�	}�;!��&[R�"�,'����.UC���I�^��t5I��^�8`�ϯ�w)���W�7�!G��a{܈cƘ[ǯ�u���,E��-Ibޫ}d��k��;�鯥��+�����bʾ���C^�]���3=}�y^����b���e�r?,�Ri��=�eT�6e��jI�XP��Բ	��v �LR�
�b�L�(f��O,Aԁ����䝞g- H-�`B72�lS/ݯ�
����߿'+zN�o���519l��E�|^�߹��5�&@�I	��Em{�
qj/Ffoe�C8�(�8W��p�+1Q~4)�������)��O��v����I�?�����1;O��o���8V4Mqf�R�#��7�q o�eB�<m�Vj'��fP��ُӬL�ۅSfo����ITz��+ƃ��,���e����r@�b�6J�Q�E*D/�0�vFR����i���m��?��|g��D>��\������ΩEU�W1��LX��̰���@=��D�I��]�b�� 3�ǐ�qF�n��.�As���1�y�y��B���9����5��=�&D��ڈ����7%�v�š`$М��[�%\�U���Ck�د�x��Dc��\������*���	g$�ً �	�h��j��F��d�W+�
�����2�Ck�)���N��%�qΙk�}c<��P)	ހķ��u�5���i2�- ]&�����J���	A���j��QqB(Y��hֲN��/�,�ޗ*�Q�����3ٝ����zF��Ye����	�vφaדg�6�3�N퉀�Z��~"\���I��i]3�����S��H=J^�p@���I�|���ͨ98;���&���9�t���*�9�?��]��XT<�	[���qH4���;%�=���s~ʂAS�q�--�#����,�HH#w�����~J�����\[ jc�@�'�2^��:j4���.>��J�dß�D��3��j��G��5 gꒄ����kx���vV��e2������No孕��f�����x[l�,�_G�.C'��p�Ġ�d?qn��'� +���hH�"��A�;��O41x�O��Q:n_����Ï���i��fI�n M���,0�T�V���>�-=q|�ENH2�������y��\�P-\K�a���'35��yd0�Ac��uIhm>����2� �|��)�C�H� ,� 4x��Z�����;�>���bm�)ܔ'�޵{E���&�2�`�;P7��P��c�80���*�z�:�X]Y E����Ψ�J��s��c��Ր9u�G��s�V������c�L2
x"޸����`�Bm�#����M���6O����}������J`Ҥ�J�z_��m�L�K�B`�B"-�G�'�b�=h��&�*{��(�F��T���(������-���=������X@��mY�<ai�t�R��V�અ�k'Jo\c���V@�C����Ӌ����ŊN�m�s\	�ҋ�"�ԟM~�+�8���e�]��Z�q��� �x{��C��j�����7l�ҜM�de�e3%�
���!��_�1I��Ď2VȌ��A��^�>s�z�����	����=�Ǩ/}=2)r�&-����M��A�iD�ܑ�vA��rkd�𪍎d))hw�=�������ð��������#�cY0�5|R
�.�|�����Ƶl�.��v7���xKb6zBqY>hX�TT�飲F�k�u�nK��}쭲��حn��[,[9��ӗ^س�j����uј���r�.��f�	�"s�U6ARmе�}6V&�k<)�ʁ(�X��T�"]�Ķٟ�����c���J�]�����!�)��&���b��"�9�Z���a9D�D9�~�i���A=-�B�W[��G�[Q$�b��U/�M��B �r �?��#`����X!�D�� ����Xg5t���v��.¹�����S�GO;�Q��WMk�h����xZ��J�䝊7��"��d��RF�\�ѾZ�څ���5���t�zӪ�9S�_,㒒	��;�R!8}4.?���"���T�u�ܟ��N9&f�>P<�?�)��ν�	������q�q��s��^ZQPM�i��zh��qv��ٔwO.�B��j�x&��_{��c����Z��)����;&�� H.[���L#;���鞰��.{��D�Dk��Ne��$�'��>�H$�S(��wT�����[Ӝb#*�Ċb�QT8�d*N����"�A1��|�A�=�t,����3����		�&V����;5�k��9s2.�*������F�6w��؟C��t���IƸ���g�u�U�����NC�lX��j?%����ِ�$T{����ɹo�w@�=���+4�AAz�Z"�=���<�Z��\�V(P'�W)雞`��[%����܊H� �G�̳\w�ɨ]���_lY��b6P//{Ӭ���OX���5�[�w�]���x���6��O�^X���$M��g.�\�,O��2s�)X�*S9����5ژ��.Mo0t�,�s��4IN���	|e|)������|��D߾�eq������=���~X��PW���x3<�(�j[q���OC��o�8��q.'g�ȏKf�jZʹ\�@�k�d5�pm��_���&[�u+���V%N�˜Z%�ދ�^�s؉k�� �i���\�xj�#^�\D@��Ld0��K��i��Cb��-?�#�h��q�tƔ�5��OM5�����@�8���ޕ���r��vZ(I���MPawj�b�Yεai�6���FwR�òNܯ����@goa�21}G�ʁ��Z��zp}��Yޞ�q�	��:»���Y�4U�Wy��AS5��t.�qho��BV�up���Z��V����$k5I!}Ǉ�m��E8,5�:r�����\C��Y{ӑ^r��TTh3�r��%�~iԇc]'F���7D��T��Z˟���{�zح$d�־(�Ò�{+�`$���.QA�O` �	b�N�����D�ɍ.|�L��?Zc�{�M���tF��H2Y����R�/C��K����|&XU��t9`|�E�.g������s�v'�L�l� �=�#�__MlV��Lͪ�ed�K��_�kʌ�p0�=up�:e���1Ԥ��W"*AJ*l~�x�xX�*j�d���wi�R�����@h$mi�Xv �bؙ����>��4�[x9ń�S��Jt�H-�u\��r�� 91`1',w\�(�حL}����zNnf�k����=���|��bԁ�Yv^�T�/=�Qq
�M�����z�	_?�S���TS0H|ǅ�V��b֣�/!�, ��Ǉ�T�
'J��LK�
�Q��C��7����&N��#�y��3��q�+ZU��1ֲd��2���l?�Y�V�=jN���h�.II���eˢ3<�}휛%���%Ǔ��g��IX�]�"���@H�* �e�_�����}�c�����=���0�53 ՔZ��)LY24ym�ߗ�P
x��*(R�\���x���/܌-�X0�Ǖ=Pr��8`��Z�l�N�����M�|h�R��1�h�(j�.����$L�6z~�
4<(CX���AϴVf փ'�m}x���"�����p�zp�!��9DZѴ%�긩��e���;���<�}�64��3\9�њ�J��g�oȠb��~X��'�d�ר	���Dvg�����A����ە�Kcyp)r�K�Bn�Ӽ��k�=�"��5�h�ɏ��vVp��n�I�z��(K�7�$���X2��($�4 V8�)EN]ϵ C����(�S�ݙ%!��m�Z�/�&�HM��	�E�q���߀w�����B��Z�{HIE�43��;.��3ikZZ�=bݟ'���q����(�����gHؤ��`��~:$a���Lw��mT8>�S��Ow�\�5���ޝU�H3Nl��c6Xl�G$�j�:y�שM��d�( ��ɿ)
���嫾e�2��^km���Z�|������}{ⱋ�*h��Y�����S#w����ӧR��˺�D,��<C��bb���}�8�~Zmx�C8g����C����E)x3}���%�X��Z����q[�-�����q����^�{|r��<K&<VD��)�oa\�h���a��u��/�*y�
Ηj���d.��t�Uz�2?<�;2�B�~9�v;�#E�����?�]�|�����޴2�5�ט�ښQB�ɕu��tޭ-v�x��>�;���ѽ�X���9G�� ��0td��KI~����ۂ�,�� ��<\a�� 5imXL�K@yЯA0 ��X�8[Ǿ����eYc��"N�j�d¶}0��v��Hܥ�6�1���K�`�5��z!>j��T�f�
�0�s���p}�VpR���~��J��Q�1-v6AF�=���\<�{ �v�½c�`@SJ��u�@�l������r��tB�gu|ĆW���^Sկ�n�\!p��`ҷ1H�G1H)���Ɋ��W"�^�'6E��y����c� �%W��>�W��u�>��XSϊ�B���P�xs����ry�y��44��B�'!%VR 	ԥ��'�P��ƺ�l��&�f�s�����Rޫ��tx� ���	��1�� �H���I��+ء�k1~�C��Η�K�J�*+.��%��$����%�R^_՘�>� ��
(� y���� d"�ذ� �j F�p����K��-6fSC����6��uҩ��T5���Ny庨�S�~Ϣ�X�d,wz�Å��Ǝ�k~��/�X�C}w'}pK)M���d}�8ǤCő�ݐ&�[��`h]Y=[��^�Y �=��T����l���;tg��ѕ�O��QhQ��=r�W/V|�AZޛRvS\��s
���L}�]�r"�>��\�tț���'-�rr@�$$���ٽ8j����Z�Km�_>c�f8�6����3Z;f����v���(����}=<!ds��^-��&f���~do��s	�����s�[��q��e��E�Mɰ�Te�EW,�߈+���nC3�O[���$>��U0�Z���-�F�V`����m!=�t#WQ��U��5�ERES8L{y����
K@f�CQ�>0|��:���̊��#��4��۝Ye�֞�4|1��]P� ���2*��{T����)��XY/��?��n̝c��)X�KԨ|��g��V��PȔ��X]�V��G�05ߊ�o�qQV���P��*=s��-�)���q~�o��C��
���t$�Zz�� r����B���[X�%kO5��I.*�p�ʏ?"G�X�6#�c�Y�/��#y�dI��x^RA��;��6&ퟹ�!�h`����xp�9���'�����Œh�����,d������.�4���҅�=.�̈́wL
��s�~�S�@CYJ]"n��Ic�zYU4�t����7��@����n�[�I��i��N{@�t?.�ay�R�z�ٺ���ʶCψ�����ލ�v�#�^��c� ^����
{��y��NS��胬}48UY~�z�e��&��=զ!7�Ǻ����mgۜM����.���%uQ(���NAKL^qb��d���H�1� ���t��_u����G|�<Ѵ1�?1,�:���j����<6l�g�p��4�(X��Yzʑ�K,۾�Z�ʶ�nB`��2��Ϙh������}ab <x$�ӾD����-�̰e�e�̹M�*6�>�:Њt���`�W���$?��%7���X#�a�kKk��-R	��c�&܍���f�h�eD����;�����i�:�F���m2m��N9d�}�W��8JqO\֬�9
��\�����
��$_�xČ0���!�=s�z_�m�����;��:Cl���8��N��D�X1騄��Qn�&�b|r�Y���L�e�I��s�l��g6��| �V�[%��e�����Ǯ�a�O�cw7R���+�A�	nIGi������d����Z�� �?��E�@4\�^�h��Q����䃝�:��]yk��ءQ�O 8�ɂ���F��p������P���(WD�V,Aa,��i����0��~$=�t�ț~+�^�H�����E|�`���*AE�9Fc��%�,X?�"8�����M�u�PZ|��<VD��/�	;�M�/:��C�|~guJ-�Y� #�t$����#����/��kO�%���\y����~4��y�8H=N����|OviٶP��gI�ݳZ�儎�4��|V�ؚ".��C�V>מ\�H����h�	ҟ�7��u^d�u�UX�-έ�Ȣ|����8��W��R��o?���0灧;�_vbQv���{X�\�2��V�}{Aڢsw���ǘyZ�������x�_�=��T�)3�V���(�ɠ{2�,)���_w�е����v.�ts���x-���6� ^�}1��Ou�!"?�<
R1�����c&A���d�y�5�vڲK��~�U�׵����3���ہ�'�u$��pZ��#n�x���=�
����1ūϝ�f�!��#��=�_��E��!�O�ɕG}����
 ���Y�Hd�L��(���$��޽��F`�+.�_S����������sވ�6;�Y��*d�dt̲#B}w�ai�z~Rt^� U6��K�^z�,�쁊����0R��󦶷�K�Rb�"��< �3C,g���TH���)��-��WO�T���\����
�(_շ>����Lo|2){oocwr��;H=]��j�����3�Ӣ/Gr����h�fr*ϋ�,;�u*ڬ��������IU�Nq�bW��*��B�J�#7���
 c"��[-M<�h0�Rܲ
�|����(F�p�5�q�#��'�c�8N��s��V=�v{������8ޮ��Gi1S,��piv�MvS��,~��ĎQ�Ԅ|���m-k�]�g�p���wt9�g�Py�(�}o�D&�����d�8�҉�<�!���|}������*�|�x�ϛ2��a���}kY�R�H�z�����&�5�Mr,���>�sn�p�r|Hk��aU����;d ���}������|�ԥ��m�ԗ�����')����Z@���7�ퟋt�As<~N�F�B��0�1��!6�{�䣄�¼$��+}��me���д�d�����EC`s"#_w�
&���&O��=`�pi�e_��(tLPH;�Z՝un�(r{��\ߌ_}H��c�[,|�>��-���j�#���%�lk�h�kd75Â�?�)�٫Y�8��ҹC�{%{�._1��I]B��fh����R}RJe�ڗ���[�m�<j^����guƛr��p��n��	֙����6��`��f��<P�	�8HW=����2E�X�g�z�˷)?N��u>�O��Y�		�p7�0ü�5�1ڢ�#0CZ8#������9�|��	��k��h��&*5�!�fJ��� �dGQ˧&l�<��u/��m��M+�I����E�Z%�(�W]rڝ��]�L3���N[#���8����0�Z@���H�0L�"�}����Y����	�·"��У�9�K���/�|�0��x>Z��^F�i��e��,���swidUݎ�v��w,�QF.z��*��tԴ
�+s��x�o94�zWʹP_~���W���E*�n#�� D�#x~�媔��S2-����2��z=7�=�h��T{�[�|_�����ۯW
���·��gZ�>�Iu\Xb$�RC�@��[td��r�T��G�������΂�5#�¥�]n�����&+ k<����l*�.x�M�w��c������"�����n����9�6�"���jy�)����������ջ�����
d�d�7SR�s�}F��[�i�c�(��`��W~��a�V�h모|\�u�KE�S_��Ay檮,��E�V��,��j��Ͼ?@�����Z䣾�����V�4]�x�Y���s��FH"���L��`�Ӿ�Ȗd�K�{E68~�GO5��V�K>�/
�H��F���;���U"
�v�J�
y *Y}�(�X\s���n�����B>�&m`��#M�))��x+����Nq >��7� cb0��i b�����M��_�v��n���"OT�|�1ڍXG�W�#��<��m�ˉ����h"�����6k�8I�39���\��f���8�AbH�>rH��`�3A���n,lД��y)�k6}B��#��o�At6�uv�.��0Hkq�E�C�@]��4� Nb-f��4C��r"(�[� =5������B���ߎ�A�ut����%�:��~\��<��i�o}��?��<�X����� v22�w���?�N樕�"��Z��	?�Y/�t�謁�#�9��ƻ9a5����� �O@�Ɔ����"�k,o�G�G#Wl��ա��'�U���ɷ���!����vcV������h�'�HV0�iLr,A.��Ë@NoH�j�x��6����2ĜavE��1Ƚ���}_�k}|�>@��أ�&?	�b�X�i��;e�/][d��!g>?�s�&��%�Ŵ��α�[��Ab�q8hdi(5O+�~q�d���FK�\�4Z��$����Xj����l�޾�X�h��k�ß��\�����rFg�ĳq�ʐ�S�����h�)-i5��
MhŁ)�ț-g�5rޯnM� �UfM��%UGձK��rA8ho��}���y��_Ψ���	�� Y�֟��g6�(�@W�O��>����s��}�6Oa��y�yW�µ� ȉp��Y���)�=]�����])*�h��aC5IK>�0G��Y�f��*l�K?y$��[7B�m.*�'?L��6J��Thƻ�X�,?5{�C�7���!���`����jz�eZ���ζ9�p�jΐ!�;xx䃭N�b}�13.��bW	4�I�D=Zq����(���}Ps�9"��xہ���v���_w,�ڏ��׈�.��E�.���p19j��1��=�b�&Q_�è�Z�6�RD���5�I'���,)&XH��0X�qKtӜ�cb�� ����W�b�->i�$Ѡ#)�̼��﵀^��,���O�ABی�y�5�]Pm,��C&����\ �د��0�d���_H8~��rz�G�+x�cDCl&���KWT��A�g���hy�?C�R�1��Q�o�|���+��9�_�:�^�@'(Ҙ�4�T(��8*�k9z �Ź�8��6k8�Ǻ�spݝ^���g.x@ѐ]*ְ;Ԣ�o��MB��e��jda�8g7w�]���/�w�,�`�NyV2\���S��ܢZ��'�aӃ1�d���L�4��2�~ǻ�:�O�G������2Wq�T5��ڷ��\U��S��zs��L�_('���Y_���^�ͨ?�wJ�G��k�I�n�����${�Q�6���;#���z{����=c�4�V�,��Y�� �Q�r�N
����KX����[�����S�z-g������ߧ����ՙǾY�<9UƯZ�M/�Áf�%�N�T��~��J��K�K\k۰ů-N=!���l�׌��?�SaW��S���.+N��R��S&��X���2�s�~�}�c�Uۙ�Z��s`��SZFl�tD/^�n�^�di��Xk���4+ө|^�ib.����]h*�����W����K���L�y@�*QSCccl���?�d������$�\�� ����4!�S�9%��TI�Y5�-�+M�⩺!�6�y�^:)�E�Y�v	ޤ`"�4��^�r2�}�r��+-��>Η=�h7�#dr��qg1�zX;�l�MM��h��yE>��{;�
`�����_2��w7�*�7Fg�X��g9T��s\�i<'��@a.:����Д�VŅL��0�`kY�d�d��Q9uc0Bk���u���T@)����iq�Y��Q�����sQ.䒕n��x#�P*ȯ�l,�-��@�tHj����(�&3A8�Q;�C��_���'��~W�HT���h��F�T�cWl��S���ߛf�X���ܧ�7u_��"�De��_�E�'�z�̒�눵���gÞ���@gl����-9��,r{`�|����.��������k !�R!���a�W=phv�c�ـLM��W;'�㇬nz��y�SUҟ�z��Qu�2�<�� m�t<%���Y\��l����/��ͽ����aR�����9M�Z��x������O��;����Vq8���^��{�
L��U:jeh�m��һ+��'h }�&�����*�-��'���M4t�*9>���w�'�"G�s�#�fhg��r�&ȨE[��w�}�&�m��/���HF�l��)H�xi���z�NxhN�n��!k�m�*�^�N2��j�^ւs���'^����ʻ`���#C����}��{$����8�̹	�	��]�ess�H�7]�c�j����0Qc�{t���h^�,�	Xa�ch[n�	�7+�=�HDRd���)Qx�w��^ �!�u�s�r\X 3�|
P���{��  v(?% 1'��}��!Q��\��њmF�j�K�Z⌼6Nm�&+��Ӛ���:�(������!��'ti���7��0�YjlK��Կ�����
��%gK���yJ9��~�ٍ�Sj]M"r���o"TAQ�ͨ�'���vSb�����ePH\���	%cU����(v�{�_�a>�}HI&V������>�XrC�T~3r�l<���C��ЈB����(�uj���c.IL«��/Rxmّ��T������X����� �m��6�X�c`J��5T����o	3�3^��b�`��~�;-�H���"��.�>���&ڗ�`�ua�V�P��&ni5a�Կ����T:�ݑk-o�_�������Q��8*�1��ay2�EM��I���	����Oe�n�\eJ�+��e�zo��Cq�}_��\�ɏ�g��Nֺ!��l����V��<�~
˕1� �FJZ�P� D0�<��7��t��/��ס��?��<C|��jC	����W��I���5���ew��}�>ut�<=5,lߤT*��(�p��=%����.�)3�yߓ>�j��&�]
Om�JU�iO~Nd���0X��?�KW~?����4��9�"��jZ�#:�DK�>��8J��ΰV�ڵ,ެ��<�R,0�/Bɥ��6kKϏ�I;VE�vgU�-���E?ULV�����(j畛0�#��} .;j�cO�ʭ�s� "ia�1�fM��M)M�ߕ���:8(����W��e{�n�u(�վ�6�w�)�}�q!4_��(*&�H,-�8d�XIU(-�	��CH�$�f�}������r��)n�z��(���'��	��0T������߾��w�RW.�*F�"[�L/�j_����]lI嫷��_G�Z��`�����DkB��V�U�Np��%ߦ��:T��\*����h��&�p	㪹w[L;gn�gp7���g����6)�s!��%�A����
�*�ػ�O�qEAu���& ����.R6UIT��[��Ρ���_��� �(���0%�٫EK�ĬU�+�"�fZ[���>ܳ}�Y6�<}PķB�U�M�cdի�����s�+:�?8Z�A^�/���M�@�w�Q�)hē) �����S����s���݈�NK��'���epQ88��j��2���c.����cvl�E�"�vD��CJ���܅�[���b)��5s������$���e<�@)B�Ր5%�(���&�w{lMd���)��5�th��R,�@��=��n��`��o .����K2|�M��Z+%QѼDc�$%�� #$����-�V�q��&3q���i�XW�N㖗T�����7��z�r�î R+�g�Q����Y��}�$�
�e��̂oTO<�K��[	=�1� C���#mo�	�(��I���'bq�&���+k�{��D�!>��s���d��7U;�rmJ��0�)�r)T�fD��_�g=�q������ 4GY�b�l_�ǍW��:����U����#n�1�%�ݞ�;IL���P�/pŌ�exM/Ps�9��(�&�S2������l\�����\�������N���;K��A����RiI�X�{�5��vj �����8;��T!:/2����e��S� ��̍(��~���pUJ����������:�S��4�1�rZ��Y>@��Ө,���b가֏�;/R����%u���)VZ}�+xp�����ET�5�g`��@��H�{Ȥ�:P<�PV��js ���oBP����IkT�^H������*����ω�nB�A��"G.Ѷ�9
m����̍�F<e�N���\�ן��aI�Bb��?���g��Ah��bw߈ H׆�G^_�h�ad|�<�;:��j=�G�3��-,��U�B|_�ޞ�o	"鮛�`U����������� }I��b��"M��CO�V�!İ��&��K3e�����5�ܶ���'d-.!�`C���j���Ciz>��@�l��k�0~�]������k�璎����w���@�uS��sir`�[竡ۖ�`m�/=���[�1���7���	d�uG�@��WOiCLL��g� tvA(.?�,'&���A�OЫU�uC��(WĞ5:%��D.87W0�݅��tL[�]��`�?g�Ӝ�C� (1Π�:1�D�G��]��Y
��*zT8��k/jNv�C����҇ڝ̛�Rx��L�!�v���a��
�2�[j�3��|�L�e����%.��l�!?�R��9K�(n)͘(ӳ%�_Iݜ�
Ff�}e�/��۸K �3�n@9���H���^���
�#y��Z,l<�Vp`�Z�JYb�����M9�&�7
,&`�ZVR�b�tٔQ��ހ_1�|ٗT�g[�����ސ���WW�y%M@n^jBJx���ř~�n� �,)�Io��y��V�>���>�t/'S�ز&�5�����	E0[˨�@e�~��u4�����X�����,A��l/�߭��1�(@=�`���R��<��L �E M	���S��7A�w�L=�pj�Y�w��]S���/q��a#�*'Rq���g�#@�J�P�| �����n�~�5O$��_��n+#9n-����k�j�f��ZV�к��=� `���i�k�?�d�C�7���7~�v!,�4��4��
� �g�ޚ�pIbi��o��.�G�}+ ��;�0Y|n���kƀ��i9�\���׆-�Rf��Г��N�0�>�Y���1H��5�ˡ|8�-(�t��O�4	T|I,R"�&l�Kg#�9��֍�/M3ҵ'���Sδ55�oOW�j�|��Qd�I��*1�Y��Z�f��<X�v� |�v��%{��`�U�;Wy*8:d]���U�_���@���"l4�h8�Wc��)a�9h� �$nv?.��+Ym����e��X�D�k8�'"
kS����H}�gl�qW)��Wb�2"qKhi^8�3�u������ v$�o�h�^TW��YTO&c�p]�eo>�ܾϺA�9jWc��{u�TZ�HS�5cޑ-n�`�8�3�~54d�`ߘ��A�p� 7����I��F$�����#B��n���&��C��q1�o/;Ȫ�O����v�<kĻ��D�z�?#�{8D0%m��C�.��!oᠮf��6�)�d?��UG���b����C,(am�%$�(�ҶΪkjj���Co�!������EE~=p��a�%������;���S彚4 @%b��<Og��'H.Z��wO�CAݻ�i�s5=$H�K�{�;Y��EU�����
�l�RK��R���4�<����|T�N%������������?�q F^��7y? ~�sW����4���suh�Em�3�������zP샥���MW��O�4�c������ˡzTvy���3���;J�JZ����v����H(]�C�u��.�������@m�Ǝu�f����]�#ݘ�{:��Ӧ�_��敟��92��͍_�;�G&����{O��{��֧��h�)ՙ�V�3D�Q�k+Վ���������F-�J����*+����M�L�pX�kn�N���T~p�� �d���.��cK�`���"�F�пn�)�;������6��*ͲȊD5���i8�ܞ)�� [8�6��Bx:3�'�h���Y�)W�ܢ��}S��=��,q�`*����Ȉ4	���O��-T��F6F��SЍ
���v�\D)���]kL�a�)��9�_BY=��V	�����b�;��zup��W��Vi�l%�C�C����#�v̵�ͣ����ɧ* 4d��	��+���5���D��!���'mL��2�-.�t<{=��h$%E�D�(D ������T�g�h����g�-+����Joi�}c�����W�7�'�W5a�I>����t�	����}�G"(d��Q�lK�~�]2�}���/�C>�g��qvq |V�����9�E����o�/�Q�J���9j@�îV�-ߞ��硁��(�Iܮk������,2��B���oⶏj�?��l|�~�Kj�b��1�GK�U��aͭ�ǒj���!
UP3gA��b:?j���\���$�����C��~�`0��Ro�cM�6?��U�h�v�&jL��m�����`N���K2����v羡ɗ����C���˼[&%N\��Aq؆Pr�x� �H��H�U������E!9� D9�Ǝj�c!�	�C֋t����;e�XI�ĸ�Ъږڻ�����@��Y�C%$
T��7�S���p�>`Hmbd��bU{��NK>G�!S�kI�d��h�T�,N�cJ��'��&��p6��W%"��a��-XX�3r܅l>:(��|RЍ�K���oz����VdW������+�h��Ʈ�Yn���b*xUƪG���V�=뼢`�/I�/�J�5e7o�1�E����O�Т�C�����������V���x�k���[<����F�H1E	x�Si�D;U=�����D��;j��e�$�8�yJ2��X��������\�'��m��� �N�l�B�I�G�p,/|6����P�y��3顝O����9�.\�GF�t�/�:�h����ç�����Vf�o~����8��
�5fA��o޵�#�ݘ��i��Fxb r���~'�9/>�kQj�F��DF���K�
���ܢH��ŷb�B�5R��kLW]���ot ��W*ҁ����,�9�{�(�%��|���=������C�/C[OƆ�[9�[dXǒ��F�)���eq����G�����#!����P��2Y�Y7>�d�T܀qx�7��d�X��ݯo� ���³C��d��J�8�G��W��Lg*�&�.�����r �����S���9��dJ�q�eil�`/�h߂�D�"v3�$�_{�e|��{0�d}N'��ܔ�b�ގJ��U*��EC
L�n��C� ��9[�z�u6���tR�e~ǯp;z�j��(?[=����N�����w����]���=��і_Gw�=�.ب��|�&�*h���R�r�E��K�ʾ����'� ���V��rhT�]�;����)��o���D{UJ���Oѷgˢ�z�t2w�Ld柛HB.�G<Hl�#@�ZY�j�hb+�P���hz�Y��g�����[���,Bk�C+T��fD�����%�T�)�E% ���cN̰V�I,烀	_}�%$�V�� 5d�"p�:Fv��U.��5c��*�p��Y����i	��"�BXz�mz\x�+���|�f�p�{"
,�E�ݲ�06|]�ոk=�_�!��P��к0 �Gz	JR$h1vt��{ً[�#Ѿp����}�Ƙ���n�"�F���B�2߃���^�OzM���1�P*����Yd�`���;S�!`��P����~���Aze1�v��!��VL��ち�-N5�v0]���c�����K�|��(QEi�u2�1�f#u>��}���bZC���C5�������P�ͫ0�]Ҕ�9'�T�@�;:�mf�|��ǜ( 4;o`1��qTJ��#��Wv�>��QG�I�[4&drO4ℯ��S�=ذ�H��vZD54��[W�c���[��*^ �e|����*��<D�\�v���y<��r�x���g@����[$��d�,����TU��ND��/U�����!i��	���Oꦹ�,no�^�H%wVC���{Nā��R�$���)����6bi���.C�$ğ���J���Oz��^2^�X1�i���v�����8�Rb�7�����ߒ�:�C��jХr�-�=�ͧ�{�q���$lk�_��ErLA��zR�0b���mX��������VL}>I�����U����`�@
������e���Ϙ~2� �򄮫gе�oG^E,G?����6�q]�v֩��	����p�V��*K@O��c������Ũj}���R�+��Vt�Y���~�h�N���G7��d�b-���~�T],�R�H
;x��6�� B²�ߗ25�G��-b�\z<�;3|���*g"��L�JtY��2�r���:���n��! 7�����F����ˀ����2;^t#�$��W��$�ġ-����m&5��Ê�dx�78�b �'�)c��m*B�Pޡ���;�/dܕ���Z,��0��٢m�7���d�y��p��t�<�#\0�s�p�⯙�9
�AhP�)SgO:��I����8*.wh�?8���L���d����ѡS���r8yX^x���E�b��G���COV!t�ΰ�Z񭁞��@�fA_KQ9ݫ��:b	����U/o�g>s��nIc��39)�|���*���|b#0���=���n�0�} Y�LњIW�=R)Rp�#;'p��}�[-���ۚ�(�z�?ި-|��&*��P��ȕ$8��Ņ��&Eq_] fć1w���(*�#�.���B- ��Ƌ��pHy��frx<�ky�*�]�y1+�^�d�e���z��?`b�ҹ�-� 1(�	��6='���\����n�4�&���D�<��׃lR��%T�����z���}(ƞ�~L�3n<(�v濈��X=���abu[����[���}�	zS7�~燷h��xd�����qW�1���DA���-w��d5e[��u��Z}���RN����vъR�7WiYͶg?���/P,���À�륖���̿���cњK@`O�\�F.^D�7�u���o^�������L���x��4��[�{Ή�-H��H$��������#8M��S������
d1�`<��Q�U#���:���Sj�����$��~{��2�8�����7C�`=���3���Wc���N�@7�J�H��������c�\��8��a�x&p|G�v�ua���.�H9�)�GL�i1��^�v��MB�ũ���/ ��F�w�hy5���-��ˊTP$�p!］�C�B���w�����4��9t��SD~��� 1k���39G������I繧V����A
�~�Z�s���e�Z��mI[oU�>v���۩�5bމ�\n~��Z,�:�|�`� �N�^�P����Q�F�W�'3��K�18�P׳߸�a�}�h4�F��+y���@�^Q�iv�0ܹ��񸿵h��'/��{6�T��7lI�I���0���5x� U���n���fV[ˌ���U��6�B��?8�&s���A�ir�%J���l<�wE\�8�yu�TO0;l�
����`R8���D�;Mc(.}�uQ�j�o�W�<��x�g�Yc�g�Ah]K^��y�咔(�J\57����C��pp~���n�*V��%�;Ԡ�&vˎ��	z�nG7j��J�����I�NS�R�ߤ�@�����B�f}��	[��'���l+��"e~�8����~�����Q�qb('Ɂ�62O
�f.��"m���JAl�%"�]��V��z��41O�U�?O NI�ӿ���}	�;E���wq��l��4���#c����x��C�)���gs��A�XIoˈg��e��R����Q)h^%f�V��ij�o)s�5RFz���Ї�4���%��B�{ֱ��B�%XS{�8���A=��̓H��� ���,=ܫ�bƲxGc�ĳ��;&9�Eb�*�2I}5^z��-Q�]c�̤����`�����吞��[g�.�i5�A��&��������ډoox����n	쬐5I!��q���J��"9�]@���	ip�{Xk��<Vܨlk���t����K��Sjh��@0O�@��$b����Ŵ?]R��}3{T'�[�� GŅժ�S����̪�^]`����OP�r�2%n�&*r5H��ܸ8���Y�H�u�����^C�������v�ab��_CG�6��K�2&2�S���l�4
FHW�2�n?_��wi3G�K\|��E/q+L�ʀ�u��F)M�J���aP*Ҳ�mG�uj��;�x]*j2�V�g�(��x���<Zwӯ��wKV�պ��r���ރ�Ը�L�������(&(%վ��Ө�P̱[f4@�EV�����asd,U�R|�rY�����h��c[�V��,���J���Q *�Xy�<4Dj�RU����×
p�MV������ ��)�e\�I% ���l�
�<��{u0�u��?�q����VH5�yݣ���o٪�i&Ǒ^I=C�N�U�u=R�l&I��ڭ��$R��φ�r���x#���8�>P�c���&�9�*Y�Lw�J�I�o�?�lR�����l�� �a��y��&�|��VG4�r2/��6�[�2�q�91yā��ݩ��:��٬���5`�S�ɣ��W�m=d���8ڕ �a�P�3HI��Z��S�E���S�$5���p�w�Y���{���F��J~���S5�˲Y���X��G��`�����f9G6���>,{&���V�1tA:1����N�ኍ�P7���UL��5��G��Ƴ	�Ntͨ��`���L�!�耳� E��[��J;�єK�R$p�+�
�/_x��a��;����]0��L���mRk�x�I�1�֨W����������
�#2��v�QW�mf4Ǝ�;�MRň�>n5�"^:l���#����Kr{t��s��pS$s�MY��<���*�*GFx�,�g�����1贴U��G(��^��0V�����P��5ve�u�~����D,����oY�-[����lF�_�[GS9ٮSw���6���A�~�O�^?��p����c��f�����_��+�*g����o}������������i)3f-�?F���-�R"�,^7L���u��z��/���Y^\��'ۡ�ڮF'K\+�-�3��v��2�j���ܐ̙7�����J���h�°9�˿!t"B}h����Z0K%2�k����-k�X���?�c�X��%�GfF����2z�a'�Զ	8��ۢp�-��e'������['*�Ѵ��^�ݙ{ΏԱ|a�[|#K�t�1��d	����[d=}���mc��B,	����U	���al��3O�(?�;�j&d��g�aֻ� ɷm���f��]^n�~���T��I[2��xA��\�������LDp�-8@�Z�DI���L�:�ԣ�*`M(O�.kp�,=$�0���G?\j5�_�������Z�j�d�!j0gC*�0��u0�U�����pw�fu��޲�W��IN��0�L�E�Z��0��)�$3�^/�vʢ�8�f���n�N�"��&&��Z�K�W����>It>W(��X�,��HL�"�����܍�>��7��ֳ�� [�6��ْ���E:�`&�
��f��T�{S�>VԵ��.�N	���ki�5�X~��&Q)���qgj�vF��eyeq#���P"@���/)�ͺ�r��I���"R_�:�!U�-]>���d������uw���U��k���6;�OK��b=D���Y�ȹ� ��������ԽJM�^g��?�2�hdx8�~-����%�}�a� v-Z��1����Ʋ�g2�g����S�Ӕ������Y9����<�kOy*����v�}�#M=>�W�-P�!�[��	��̵�
��l�% ��(��R6Y�t����^
�ԑ��
�@ʼq\P�rȚ0w|��/Y}0��P<���t��q�6��u�	�P�m|�`]�$����q>��>��J����2�.�it�N�<�ͺ����Ru�v�+O��o7+Ԭ��	���������7�sq���r��������D���T��)�-��j\����?��5C���p�k9㉣��-���9��X񖊭O����D�pG��û3���ـP�����xB���Kj[�M���e�V}��6`�!%����35�,q^4k#�R�@p[m�A<�g�d�a�H��[x宠�JV�$������3�ξ�HMH���m����F��瓳�q̤ =�6����b�� ��N't��'���`�֝��2����m���?:�t3{��({З�����xl9>�s�X����7
���P�$F�,�j�)LyBAf
pFΈ���"{����(�S���K�XN�������`����0���؁�|⪵{6�Ŏ���PY�� BA��I���X?��7[�!Qz�Gޣ�ĭC]��ܹ(�Lw�v�������B����{��K
�"|J~bHK�E$�e'i�y��/1�.��G�����>&6=Ο.<�k�a#�)E,�#ߎEk�0�C/n[��p��|x3���F{ v:� �H�@z������D i��_����}4��C�S�R
:C8K�QZD.�/6gz+�U�n ��%�M�_�� 2F��֍n���0
��=�y��N�\�������S�����%Ts�w�����y@=�/��w������kc��~AA}���~̝ѫ����ܑb��N���ng�hI��^?.�f�D��.��3�0�o���E#oU������;,#�!I�Um�l~ �� H�nT�%����� ��v�����Y��M� E7��2�)ӭg@`Ejf%i���n�Yz_ޅ��0�)��[n5�Txlf��|�wsS��������*l k���?���J��8~�cI�lPJ]�����V�2!-�=�3+\"OP��;r��W�;��@��G��o���0p!9��jY1o�v� t����_Io�����R�aZ��<w��q�)��,i��z�T�Z[0��Q�����Y�D��-����'��W����9O*a����p���'��D&e7�����S�:��܂6g��o�m���
ѱ��3��A�c@�=�\��6�fD���?wݿp�,-�x>��]>��ȷ���w�g���]�:�g�}��_
b� �>F�\�]xe3��7\ƌB�k��4�yZ����?�͐�oI���!9c�c(���L��$�;�-��D@\��t��T�@����5w��'�`U�36G_�ͅa[���J���.�	�s������;v�����pʗ��q�F ~���LA��町Ȱ���/jLd"�Q����1�d��D��y7#	���b��R7������F����)W;��Y��:�;�,�6��^�E�M���0/�4�ǡ�.ȫ{���_(h܀8>G���[�6
�ۘ�#��D`�3J���Cܲj7�7�.6��n���~��`�?�)���*��k�^�s��+F�y�L�vsS���N�^��6/��uH4\��-޾"ݏ0��_�V�k�jd�'-��QvsK���7+��1R?��9gt��p��4�ij#/����2���~��[/]Z�/��[��$m�wu-_�/W���L��{$_W�D�p���?U��V"T���,<�,�M%J�|9��iG���ى�v���x���/�A�8���_Î���U �5hpf��`8<.�Ts�	n�&��QҮi+�o���]�^��(v5�,�g�(�k�ZU��F%HW�i�v�+s�	���`�b]�ꎯ 	�|���V~1:�Н���cY*�ۈ�{Ш�mN�<��$h��>� h�t�I�Ĥ�=�	U�i��z.�Yj�zK2����x���]y�!\o��j��ڋAC�+�M�\�W�p��Eq-*���K8�4�l���W�12�.�c��F�1�몏���u���-��=��`��*�g��P Gj+���,��_Y��� �)s2Z1�*+�8�h̖�i�W�>w��}��u��C����'T���E�F/r�������-S&fp�P�|���-DE�;YOQ\܏��ܓK &�%����T�� ^Ӧ��h�n&�:���Cod>Aj�g�ߕHI#���b���2�Ϋ]�Sq��K}p��gj|=�HT\<���n��^n?�&����㞑�:S���∛�:�\0��x?p�J)����|�E���}0���[*�h��II��@ć��+�k�̅�c�:�����Y�/��&����v�$ץ��@g���v�x�.��@E�͵�.�PW�ow]'ɖT�IY	�c�����$t�����������I}�����R9H< �«.�ZDׯ�u���i�O�KZ�)w6)�JBL��a����0�΅G��"y��6IX�&c��,�2���l�z�_�6���s
�Duۏs=�`9_��S���	Vq�#��NӦqB��mǐb�6�D.��QHk�R�LFB�c7�+�f��.��z�L�~Mt-�3��D6B��^��0�#�\�I���Kgu0���Φ �pĈ�E��N}��1C������k�x�3�c��&&/b�T(q�g��� ���I��㭄=jV�t�Q�d�D;6B�U�|@����UW!(L��{�-�80d ����t�yZ -Lў�	�de��������q�/|a���2n�!?=��	Ee�hY?��qV1����kO�I�BY��Z���,F+$��]�^B�Mbρ��v/t\��'@xw�at32��@W�B�GhG�Njǔl;LF=����x9�����ߛ:c;��7S15�bC5�1(��K:܊�e���6]����]��y>�����6	�!ͩ)�/
pHk�t��{�K��7�A��Յ�1RO`�H�K!މh�Q5�u~Ί�t;J��&e��1�N֓�~�)���N����XE���)躠���v�U��~�����G-���� }[��U�l3�?�ޛXc��(Th{�$�_�>$v���7N}�=E�/ԕ��b�/M��ɺ��Z}�ƨW�bS�j�G'f�bxd���(�`#&%o,����䚡����[Fx0�-�n����XGδ�dg�p}�ǩEt��*��9�T����٨%�Z$X��\E�
/޷�Z��;����L)T)���y\Ҁ��[��� �<J�k�ڎ��<dv��k��\�tA����=���.]���%�I�gw�G83̘&�Q$��j���&랛����*�S�<���"Y����Z�G�P����6:���c{Ӻ�&�߅�O� j<)�A�l�0�}g&��\�t��GC\������w�"�\q'e�_N��K�!G�}Y�۴3�WǺ�0S]�Ԁo&l��Ԕw�{p4���I:����7���V,= ��+}l|�_���v�D���,	��c���,/T���͇C��Q��c�*�0g�c��V�x�䘍�A�w���3��G��J@����^oz@�642]yj#���$�O�7�����A�qO9�kr���� ��qT�.l}9��wa�P�S�����#�:7Ţj��:�)Zȶ_E�����N���1�BI Ō�s�_�'U�sƇ��e��s�L��E��S��佖"كZ�0�>Nin ��^wK���^qF�U�$Ug�-���y�������4��� �R�z/�p[x��]NEQ7e���n0��L���r����P�����M$C�~�1tX� �Q������EG`Y��=R`_�cFfg��Y�fuI�=����H�[pf=����O�\%��v\
b�ik��b�fKm�y��X
�G��~Ȍ�J����a
h�U�$L<ҽ_�w%-�h���⎗�^��˴Aܐ�oEq��ZH���9���3%��N^�sk)�=H��W (��/Մ�3 R���"���I�����E���,�	���&5Z!���-��J�T��D�j5X����p����;a�P��kxo ���|�@$5ж �FN��<�nW>LjG�g*�_+5f*iQP���'8�n
�Xm���HL��?>�"�m�"*�e�Ф<�[x�^d��i�p�{����m���g5,��~�#��E*���=�ҩ#2��;X���q�ˤ����v;ِn-�Ht�3��M>i��vaiѭ�#�*U��HⳒg���Fw`80p��]R_�o��?떡K�mvW�J�0��SI����iK��{9�_:5{$
�ȕպ�}'�}l�8U��k.�P��+8?�����VJ�������jg��|����P�qq�|8a�Ͻ���Q��6������/�����:��J����;[CK�zyj��G�t�$e']f�_u �(�d�I=4�m���,������)��-S���e���t�bXr��{�5��!�Y�$'�[�'"���s!53MH �M���mKZ[.��0���-��Sb�X��O��/�~f"�ds��B���c�b�������֗�vP���	�g�o�
sx�\� �{�-l�s�B49��`�^�i�PL%o�O+7C#6��G���8���ϣo\̣�7���e8�
���5�r�o���`Pbw���⦫���'��R����,dL��;!X��Q�{b	�l�i�L��v��g3��T�Hh�^0�{.�m�k��e�6��\���%/<��@��u��)��]�
���y5t|�����J�k�Y�� c�r���e�N���  ��Pa�X���A�����8���T�U+���%�̓��e�S�����/=��I�\�����@�.�<y�ρo���	��ZI�Y��}��#�8��]#S��>9�q��)�Ѱ���U+�H�H�`�m��uXj���TۖЋm����CpwVmJ�L�!7M�INwZ�M�!F�r�M	Sԩ{N��2�"�� y�Z�"�|�߯�:�/!��	a���`*��P��؏u���J���!/&Ϊ�<@��'��.v��[y��Q��R�r�xH�����'��� ���7��b�l������i�l�/�/���h�s"��7�`�w����\����B������V�yX�t��>f��i��+��d/�MG�+�[����M��:`��AV�v4�*o>�����:>�a���񅄏x_]�t���:�����aq�0^�g��*!���څ)Rq�h	H�'_JI�P��-`a�V���L�$Y���9@P����L&��F\~�d"��B���@�^�7m�w���0���7x���z������/<����;<� g��N���#E]�6Q���{d˗��%��6��m����[�8Ac�N�.�D�l0��PB�˅�Ǝc_�?��z���3'tM~
~��1��&�oa�/g҅�t��м�|��R��z6R�ِ���̱���:#��ļp�$U��[(��N�+���|(w����k@t��㓢.Zs�ԻA# Ct~�|���e�oJ�M4����� ��^��>EI�xʍ�fͿ�}�OY�g�0I:�	��]�ӯ�A(D�kr�.p�Bүؽ�{��3Df��DmiQp�4�18��CQ��8�0�eyczs�={��К���"����Y�n�����A-���"�la�뷧� �\\H��[`k��𰛨x?S��,�/�L�'�NEu���ڍ弌��#z�q���k�,�z1m	p�E}��~�)�1���u��u���7 �%a��^b
�I.���ɝ������$�������j����0�R���G(J���6���w�0�x/V7��(ƱN ��g5�0�0�=�[��Y.Z�Ȗjo��pBB�~]޹0f�tD ^��×�t�����uSO�ښ�8� @fPl�M��l���.������#Rq+B.��<	b㿿�<N9�����I'���^�A[�YJ�^;��x̥F9�~��ϿUH5�hTΙ9cރh2Aj������!�#h�y�?�.�m$��c�|�Q�?f�hg~������N�!�ھC�4� ��*wX�19e�����~2.%��@���9�y�z�O/�
?�䃆�8?��L��bգ���
����Tq����t`HB��a$Ti�$p;㰠�y�:~��A�}$�M���;PI��-&;%��Q�݅ǥW�u�5�\�I��Q�T�F6��i|I�`x�*c��+P=�
�;K��+���2O<�����2��o� R�e��<L��/U���q[�2��'��%�rz*$Q�v{��o�d}�=ސj��o-$>�x�>Y����a��n�l5�!���	1YZ���c�T�ۀ�QJӮ��X��ph2�� ��/���5X����Z/�yI��i�.T�U�fl:�Q���=c��j� {�Vs� �8g��Ҋ�Q�ӌ����6��*��#���D�u�YK��j�}ôv��,'�a�M|K�WK���o�*��(�B�E�%Sң���9n���Y�ү�C����2�o�5I<����3������t��͋5
��I���H�C���/y~	��#�ͼE��NZ�e#kY�B9��X��UHb���;�UkJs� z�/iDg�LPf������i���j��}<Pxr{n���/nد�G�'��Y6pW���v~	���k�?��,���蘒��Vxu.�'������$#�]^V��Dk��)�po��.l�S��R]LE�YcK��6�	���L�)d+587��������m(�3�f���i#ɾ����vO+j�eI�-F���>$�(D`�u�C[���c�Z
"]��sTAE2nB��-2�;T�ށ���Ԉy��>C0���MV��&uwb�㘕XnQW��C��W.��p��d\ ��m"�nu�>�s��RAQX�BY���<��І�x�,�v2�!��NZ�W�.0n��.]�>�=��(٢G�o�	Q�I,	!���=uې4�wO�J:���3�?��QP6Y��=��˻���p1����4�XAv�%�����΃�s���>���ڂo�b�-U�8��*����Y�(>�Qu0{���gS9��wn�e5U��������,Tƙ���~��~����\����0�jk)7D5�(@{tѶ^�;2t{	Q��l��CVg
Wlq������Fo��.?�D�\�'�ECPD�8e���Q�a�?�T�I��䫪��\��S8�G��VR��Zu��J�}�����X�'C���V�;d8�G ���ў6>��s����B��ݘ�����A��o��Tv$�� �ō&`Ls	�NnʤM�_ ���1;4��F�p����y�	rp"��Rqk�u�۳�e�P��x?-�JC��So���`�E�s��.�-��=х�3�qTྐs:�C�7r��� I���G�E��͏V;^�g�x��
���Gl�'k9����'y?_�W�`����j�_��PDc)�����B��oMc�W!�)XS(��e����c��*4���Am�`��o���*2Y�k�WI />DN0W�p���r�Nğ_[����(=�lRTu���ͮ8��R�⒖�u�z!A,+ꦫ�Oi�� @�s�2�b&���>��4� �~ե��W�i���'y����=��I��@�#���7��d��l��O?vK�mE꣺�z"�"��R�A�m�3�����'��&�S�3p?@M����7&�5Z�p����`��������C��������x@�je
	�\/�A��ܹ��HH=��Uӱ��es!Fl7���@�t�����#�;<�!kf��M��X�f����c�v�!���ڌz�	�_���~p�'��y�)a�'��-�����ht��0E��o*;N=�J��?`��=�]�.nη��pP�ڼ��PLo���ju��{��I���9�� �#B�n�@I��7�s�%�6ȅ�{����ФI^{�*�ԳzVG8�h�0�}<�Y�wo'-�%��:�єᅼ�1b@^�Pӿ�����V��yYa��7j��F?��W�c����TñH ��� �)�р���Om=��X����e1����t��~���QN��*�Íl\��Ϻ�W+[3`lJ��C�@�(���Ѳmt%\l�Ё71�͎���ֵeW͂+��?i�+6��Fَ�:{Gl�DpC�,Zt�:���Ϡ�Rz�}f�6Ɩ�5T���K+5�ׅ�WV�D�/����3��F����}ݎW�5�Ô#�����kyu�qX�	/.8;�Ok��f��Q�4xq�J�����s�e>9�rھ6�/�u��ա�HVX+̦8t�%������@񴊔���ˤ<0�&�����
�.S"'Ҡ]ǜȣ��}�e|%£҇k��ޢ��C��Ee�֨��.������~�S<j�4������u y��aK��(|�E�aAc2	��L:͡��|��>�KU��h�6$�Ga����Gj�)6��.Y�pV)�\o=kT�b� �����-���WJ����ڤ���I�����zmgjȲ�)vQ{z����j���31���t	�+j��y�y�}ab�C�f�g�U{�3	�"��9�Q�Ӄ��F�f�����#��<vA��+\�}>�a������� ޔ���cx�~5U���wu�RΨV�����'���ܨ|棆�@î�7x;.���6���Z����+"Ta��J)*�Ou)�U�kZ�q1z�'�ɵ�[��$�lq���tߐ���G�X�����T3��uå����=���0����:&�<��d��@��nA��)�F�b��2J#U�]���¡�j�-�\��U�_U�s�0���:h����'��7� S(ϏY!�g���h_���|�s�"p�MФF�����aY�S��i����f�{*������?�"[C�pcuJ�S\� D�㥶bm�<�.O'n3�[��,+a�~�aW������n����#�8��/Mw�G���**[���م�;9;�"	PY�jW�-�q�>�느d1�����O(�W����!���j��)��/��Z�̠���`S��	(@?�����C�n��3�P���ۉD���0{�:�B���k�%G��̕o\�m3t���|��6v Ǐ�$������+]"���P��+�mo��D:1&ĕd.x�p/C�<#g����{��\v��$�-�����x,;�1o´l��T��?ƃ��-Gaߡ�x�c���
^�e5W���#-1C�Jz�d넄�j� �M4�c"�:+�@'&r�~b�E2���L�>�S�2A��MBQ��$�(X)&�;���:IB
Q�����D|�d/�d�p
n�N�1��l���Y@�/
.?ϖ��eS�O���y �i���dVM�:�\�8���8�-��Z���%٭gJw���@��I3��a�����#:=�d�ё�6���o%�!�RP~��O�"х	+w��c�����X�M��m�|ØT�4��Q��RYG�9� E9�x���~}�,�^YeED���&�N���룇�G��6��0=���YZk��ږ�h�7�AOl�� y"OaQ���7|ϙ�m�-tc�^I��EB��b��.H�p��w�2	̴�$ ���z�}�;4#�#}5�h�""�ږ�gb,i-�5T�*b{�r�f�v�=]��$h�ǟ������S��c#��'�L��ç����Z�f�*pl
����d�;�,��c�7|���"���G,~f>B��0
b ��E�֙5� 1Hrg>��y�Y�h3�En�N�Lt�$q z����H���@����<�-x�G �F��ư�������=��{�TkM9`j���W|���,� �D��.}�+gG�v�b��~6[�A�r�2�����eSE)x����v�!�SI&�9���t�=6"?�D�(���,���3CL��F���"��/Y2�����g�����fI�(������X'�x�2���#1ږ��{p}�8�MNmN&?*�FR<�4,����NSdf|�������q�ݰ��pC���_�w˺��B[e��ꐾi�Vc�� c��CE3@e=�E�P�Aí|f�O1,�8���6�:���R�%��9v�,x�R1�MW����g��UK	��l���R�[)��S$2��_�m���Z�!^ƥ,�6Xz_vV_9H7l�����~l��Ǫ�����؋�oPC�%`k�Ă3>�ܘ�R�������J������m��$ojqp��c���8Al�B"��Y
h�R=e9e�T���ƍH�+�g=}�ߙ����PD��WZT����\4(�u8_������騆�4�H���ܢ �<e�@�A�&�ο!���A��9 �*a�ja�}��.d��N,�R���p2-�	�M�9VK��y��ˌ���`�)	7����8�� ����o�5�_���O҄V~k�x���f��=
@H������]<��
�cQ~!;��_�`��OĘ=3p��x������'������S��a�b,�3y���q�?�z��l�y����{ $V����/ֻ��b��Vt[������ }��.\?��B�5��9�.G뤭�,<nS$^qTyȧU?��n8����ـ��H����\^�پ���q�b�5���N�<E��Z��x���#6��T���T�X ~�?�s��0?��Cr�l��>��?�D�i���}`��<�ȱάV�ء3<�]��PٻP�V���fWt'FU� ���e�7`��#U8D����74ie�g��%�DG��&��n����T�c�U�+C��!l�|ꦣ,�;H/���ʛo AN�S�a�2�������u��x�t���haӠ����"����C�e�2�@w{���&W����^.عhs��ى|��Hc�r�*I�j��}%��@�`C�[�-4'�G#(}�4�C��5tbxF��߆
�c��fㇺO���N��>p�M�7���[|���q��H\���WѢMD�(��?���)��&�i��i�H(�]����P��zП;{-��
ZHY ���Me�z�j��-A\t	&���8���|���cR����������~���3z$
��i�}[d��̑xާE��!��psO��H?�Tc<<0��ϻIڻ}�`���g�d�و<��0n�/9���'�h�j]@��L^�I)��?6�A�wke��bfz$�{�Nwv�7��M^JW5���^��o#�h{lg���`L�]�!X�&�	�eU�3x��c=e��#s鴏hgeu����ahC����1hK�_�f048��7I���Z8�����E��A���g00�߈��$�yiE&�/�a��l�Ap��`��;������/ON�[�R���;��&!Rᔁ^�g�1ɬ-5��a���߶<��H\�z�	�'��ɛS�XnK�om������å�W�_�?�� ?j��f]�0`B�~9�: �&���G8�9c�5B�B�M�U�R'���C���	�	�)yL#fiss���7�
c.�J�sY%7|FAr_Y?SWq�Q��(�j�5�Pd��unZ�(��B�*q7�2lkWG�r�M�?��8U��IZ�~�|$ub7�x⣅+��L�*�[5�>�-����_��AE���v�}�K.K�f��ж�#Hҥ�n����d��U��,	S�bͩ���؍e��o6���[��ȫ9��#18*zŁ�Sf.C����H�G���g�r�:�n�n��k�4ۤ-��}^$���������4 6H{Y���Q��G|j��j�}J����U6�!��t�W�}�!fb�/�'�.�������`��t*�:�(D��]<��c���t���\�eMdO��:���_M��jh�v�;��,埈ƒm�e�g�R���T����E�	��Q�q$޳��2� ��*�;�^��
z�"'�����p��"N���X�"L�U"�"~�^j�jF�>�u���xL;yq��m��C��g�+����?�z|@�q�{�{y�iT�/�1:pa[Y���#j��Ij���%��Sٽ��I�|��o��ӂM�	=�����5��.j�Ô������P�hjK�����GE������S��ֈB��,J�iԚ
%+Ilq��o�� +</�j��$�S�	c]4B�[������Y/͙n�`U��g��$�]���»�-�{ҳC��D�Q�2�i=SR(11�´K����U��$F��_'�W%�ĨM��zGteS]7V��:q��tT3<�\�=�2꽷�92(~_|�A2)"=��Fo��?�]�e|!�q���9~�>� Wi1��³�ߠ�ϱ���˾�n��n�?�.�-��=���M�KbP��o���"�7�5�r7w}�n��r�\������lfYU~��QvLv�:Y��+�3�[��]�{t�R?�b6�'�x���}�u���1�%|���K-	aQ��.�g����aj�R-���S`*)iNb��ԅMl,5R�a�X_yq?|Z��J�A�]�є�y,�P;�wʜ�P2��R$\���[yɠ2��Ķ`�O�~R��MO�~�E7gx�۟�Sх�jk4�hY�5�����
ȵ)����_6����8�o��Oѡ���>L^(��:�ġ2�u���Xe��o�̸O��d�3p1o�(�=��슼S7�Ű	��~i����=�'�H�k�a�iv��8҉f�����CٸM�|)�!g���GA!�77oy��>L���c��R6v���s�ԙ�����^t�C`ap�o���T_���G�n��%�ae���տ��\*��i+�0�<1�}]}m:8��~�WW��T��~Q��i��ʯ�l�O��""#	��p"�_�_9���'o`��y��1!/�������E�<�#�)I�T�����'Κ�M�;N(*�N8�S�B"��%��u�N�O��&�ُ���I���� �9&��p)��{�k΅��g~��N�B��¸vdY�#��ޱ��Q�+�A��C��a?�� /���0i����Th$r������AO��݅E�/ț�D����pr3q0.B�7#����c��>#qf�SdNϮEk�~n뇱�l�n�7��8�&�Kl����Xݢ�/ȿ�.�c������-x���V�q~U� ;�`��GrچvA��Ĝ�.��Q��*����V-(	�Lj�X�Ƈ������Yˀ���N�����N�[&t���'���m0P����3�����m�#˕�_=[)Cjh�P�6Ђ��z��pqb�	ó��#x|��g�P���b@����YY�(�y�iy��*jo��)��Nɧ�S�)��i���$A��v^�<JaA�B�k�Y����X���*��$�,�PW�&��7. XS��&��o)���H��H:�����z�;8oStU(MKΕݸ���+L�D�Zn����L�^�pR;�ma��k=n�@�[D���\v�(� ��u~p��Y��p.s!"��nAgv�a0PkI��|<!Ԣ����E֊{����#�%�2ȭƁ�b���^{���Tr�Gz�JQ(*�a�ܟ���`h^�o�'GT	���Tt�H�oF����^�<�0�:I ���7V)]������~��=N&@�ޒ�}-��H����w�tL�뤜���?s{K���	�ѥ��f<P��!�A�9�#���ڄj_��&�dM�	�h\�3�+䖃?�bO��H�oZ��]4l>���UBj�ev���c��tY�|:��X���+<R�|��/�t�㧶0{kI������Z,���J��@�t$��Y)�}���d�(�Lt΁{��Vr����l��0��j�����Ȣໆ�gUl���[_�wa����*N8Ԣ�Wک���(���[S~������
A
c�,R�O��7���;&b��AEz��#B�C/����!q�=h#�-�&T���/+��g+���^�4x^N{���r*��(p��H���{Qp\'�	ژB�K&�n�S�Z��մ,��Z��I�W�����k�V���E3a�Pi��g��	��_��}a�ehӄ\�xJ��ި��a�nix��B6��>Cs��̠�C��~k�?A���δ���zγU�-���|}�@��|ݖE�p)�L6����	&��-y>0"��kOG����:�~�R@�g�}�b���ٻ�ۏBo^��!_*~M��0,8��%OH�ג�+���9vt�ژ�i�QW��B�+(K����o �_�
?2,�j�O9�ֿP���˪֙��^�zj��j�%t,���,�TQD5O���_]�
�~0����r6J�/+:���i(�:��y�gvvT�:VHg1�x��e�3��p�8�&D�@R�u����������iZ�S���U����~x�X.3�����:a��������m^�6j��8?G&�1YK�-�Ǚ��f��h�p��d�q&�	��G$�3n��e� {5exH�"1� ����ey�����)vӸ$2x���X&Z2�}��FU��T����jk�(�n�$��
!�!CY����.F_:�$�G;��]v^5 �d?���kd7�5�}�g}p���U	��0<�K��M���p���R�U��r/�ш��wX��VpSʌ"��&k�Xi�j�a���x�-�
��n��,I`̾��^F�f���VU�62��F�Ua�hX.�����]ȴa'�dF47��w��:5�V��=�&w�2��w��W���֏�\^��+����5G6�D�*��YGࣥ�����5�k$%{�O����peޏ��H�)��]�)�B���Xq�
��ת5�	�K�N!嬑��������>�J�ѷ7_�i��φy�4��A���������ݗ&R3�Q�Q�Ip�;�j��BWvٔq =��@��J�n8e���@���=r��������AJ���L���Y$�Z���T�j��I�Ɩ�֩�׌�sG.B*%;j�I�L;N��T��[���6R%{u'ld�(����Y�m�u�|����`|^4��k�ψ�r_�aa>n����tIҦ���~a�'�;Pkpny��#*���8��JԬ��e�b5ܾe�����e8(ɯI���0����S�u}����S����>-��c�T��q�������B�N���(TI֮	��O��:�8Ă������w��
��x��è�r��8ݛ�rҕ�A�Z�cB�L��'�����_��!g��T��C��u}��$XG���=R���8��7,�FioQ	f>N���EO�6	Q���iuQ}6��^�'M��{ˁ���g�6�����������b����c�> �s���3,��/l�5v�~�[���kw���W��'�W��;TJb�_��s�}�&?,rBm�2ɫ��f�����@,�>-�-�K�<Ww#�{�U�T��f�D���{�&09����h�"�9��K�d��6��k��ek�������W��#f�A�<5^BZ�\��i��-���`�fM��6[���/C{潗�����]����A�l���
!�Э$Y�E�"nl����w/T���j���k��Q��nj֬�|��ŵ�,wҫ}J�"�7��HLx5��Pe6+Y�L��:����P�f)_�%� H<謢 ����4#`������P�I"�-����O���/�c�):G�M"��+����s�ɽ�kH2�LT�d�Nq�Y0�p�WX�ڝ�J���A^)�U5���O1� o ���;X��Q��wꘙ �d�3��ƻ4�L�/��Q�|�V��SG[��i�ߏ�}�6�(pS:L�4�^�V'��6�7r"Ol}7�}T��-�[y#~�1{OX8�#��P_��{�\����4m�9΁y_��D��pɣF"E�IL0+sp��Z��/~��~�f�*�2��@���y�.'��4 y�[M��%:��pG���C�&>�נ=������%3�vAթ#�J��?^wߨ��ٯ��"��U���4ajC4�ėx�c�e���� u��}I�h�0�Ú��� ��j��>x�jlZab�5���z�L��<�*n���΅	玪�g�����K�1�n�����#2���Гf��.4�"�����q�:�>�!�<N�,Ro���3�F�d�`7�z�Z������IsMڋp��8���r�,��,�=(o�t���8�/="��L�34��pF��{��ۛ�4g^Һ����c����o����W���lۇBA	���)�Q��Q!k��Q?\}��-ILD>���Cz>�����>�)�a`���+��zm�f�z.�r2�;��э�u��&j���[����w@/�Y�C&�eN��)՜)�,3�ǈnw`�2:j��lT[6��k*�N.5�76�`��K�,3s!-�o�fҸ36�\�����8[lV؄����9w�Y)��D���l���郷����`ô�&R�P��Y>�Y�9,�i���փ��ѭ��U��a��ԨP��2>A�=63o ���7�s7*��w�<f�AE�QZ�~\9~��\2�Д �K'��㧁�n;����ũS�Z��k�4��p��=$����*^>� IRY�85��Md�lq��B6��u��NOߨ�eܗ5T��������١�,��v�V�d����vB�	������`Y{	�
�X��/~I��{�'�k�v�J�����2M��a����.��H�*J��o���iC�5�ӶK^],"V���u@#'��]�һC� 
��l����=�yB��*@�z[~F��W�Ųx��kL��C��ܡ�rB�!�2<�e)�%�y�=Bʵ��������>���l�:T��]	�S3U���$�`����If����� ZN����9��t���	��6�^S��T�c�s��_�M>z�6���uNqD�)9e�WS��%��2a Gi!�> '��0ݩ�[�����gN����f���a:�:1H����Ӳ��I9 Ģ�9j)VL	��������0��+�h�M�ɛ�UN�A���	�Q]6>�^a��u���tK�N$�);rc*hjwEc'C���ڳ�ȃI��. o,�j����\۪��쓫� ��Ԭ�P�o�B��c \��P��T��X��g�P\�?{L��+��I��;�h�x���m��*3����
���q�aM:\i��T̕F���gM옆!��E�nG2�y�Lh�ᨣav�I���;!�2��)R��׏���"6kl]�/~q�n�帜Β�Xz�"����S�!VK��C�4t�|"��$�x|O�}O~�}J���h0�O�����f��S�_ӯ�'ݔ[���/�j*S%��I��)������C;�:'���-��^�<O��+���%���|v��2}M�/'/�n����̞���/�pa)�����F�O�;�`@�,�l�sH2:ϖK;���ҥ߾$rz�{h���J��S�v�kfgݔp�J�\�ϯn��� �A܏Qi*â��8*�����l�O/�<U#ɳY��uN[+D�TGʥFtW�~(^U��.�\Z�����^p8��M��h�Kjo{ٗu��
��ix@�r�r���IL�\��/ܡ��B�qO+%�Y�8jo������������gWzz7��`����;.�_ɓ]lӒ[�Y=.T}ܭ�S�� �uȽϳN}���p�'��K�6�ƍ��!����N�{�B��3�Byv���F�'mCL��#��SY�L�p��$WQV��p|���cz��Y0�q>u�������m�Ll�?���{W#����Y`iH0&�����]r(PyV8X�I1X"��� %&U��'@w�a��A��7��@�{f�-36�OÝF�1�=sA{#+��Ŀ�ű�E��}J��>K���!g=�2�ZG�!��;?�Ҍ����j.b�[�]��ֻv�o�GD���Hnٺ�ȹ��C���[�x����S��+���y�����̛�l{Ţ�τڞ��� �λ������L[�����`�63�kTMS�B��'a�[���_�����͡)��?���`*z�h��`pB �g��P��LBl���v��7�Y���~��٬puk+P�솂��2�S�����[,7��h�"�������^���Z��&�q#af�#�D�=6��i�k�W��$�v��]�pU;�9����I	ڂ\u�B�N��ZO��$�E�_�{ϴ����"�K%i���t�����M<Q�6��w�Fb����l��:�Y-?�ؼ��%s,cr
9��k>�"_
ʕ�t3��Vj�� Z��0���[�j�:]��[��v���j1�7�̚��	y�����s�����wx���/�\x�F��|7hN<b�ߎ-$2��G���;��U���#D���k��o�Z7e��H�WB����jVz�G�4W~���Y]�������w�r��-5�q�V�B��@�#�yQ�k�z�������c�*w��z�����2#FL�QR\�i&*_�= �.VG��8a��E@ר��GǇ�9Ȩ�n�5�жV��g��@���
���A��Ľ"��:r��o�$F���+V|12@��l]PM���`΃v���ё�r�⺱�z�Q�)0gӗ7L��~��dyJn���M������%򘿊ǝ��==�d�r5�)�lM��M���ߪ�����,;2���Ι���cԗ= t#ʹY.��J�������󬞡�m� �_�[���,oǛ�]��R�Z���~F׳����o{x����FG6�a�Ey�@�T?�}�Jai%X��P��׊׶�ES���3+=f�z�`s�T$Q?&Wkv��񘰘�N��r8$���{�{xxi;��� eLc�ĴWŕ#�Ѫ�;��4��8���6�ш��xH٥"`	������֒K�� raN����y>�e̢�y�w5�n�i!��\hq�m�� Rb��hra*(ˆ'�(��|�C�q7�K-��ĘKF�N[D�*�|<���1q����չ�#5�BV�����𸼷ø�b.
��W�!�R溣Oe_ܬ�U�kU�� ;ë��1�����U
�X9�sE�gJ�Ȫ?R;!D(�<]�\�U|�b:�����m�vw��M+��'���1���l��B�
����İ9���U�հ*7�f�9�Ɣ�����ٮ��T��v)6ӢщJ�i7_���ZĽne�>��U$2N�&��s
a��=�(�x�;p�o�<!��B��*9��h�/�-�� N@?��GdV�V��t�C�'Ҧ�3�2��Ma�I������%d@H/�-tz�;����l��+�"�w>������6HT��iHhq*�uzK�E�Ѡ���p������[��k�J�>�~|9ރpes���U9B��a1��aM:��%#O,6��{R�����V�
ݯ���wz��>n��"э�E�dw�N��鐴R�f���x81;�1r��]Þ1 �'{\p�hkj�����$�+mE��-&Vl��O�YA���GP%o�c��%�J\j1/�R��y���U�σt�q��`���odj�d#��٩��K��A���|����+�7���aN�+ΐa��Xs�Q�L�D�z�y��x� |}_�4J#��=H��T҈�S�K�#����g��g��/�%اFʅ	�I_	v��2���ʅ��`�0�m�����<5L}D)1��D�Rkh��i	
	�m ����f��ʄ�@2C�٦�_����� S������u�wa;<�9HF.Bܥ�j�tІ�2����"O��ޖ�q�Ho�w��r���IZFaw����j���jy�T{m��($�c;�+8�t��I�5���5�gy��ƑA_F�~��pAIX�ND������`�:���� �b���e0����G=��Vv��; ���Zy6"
��t3*iJ�QY��rb�E�6ŷ]�h:��ڒ�B� Ƹ\@����W�|e�Oۢ��Ym出�����X�#Qc�� �?�'�뛞��f���h;�ac��̯�����LGQL(-�a�.���,{�pZ��mk��[���<v)��
���?g��F�����l��X�|��.d���4Q��@"_�˕����y=M�ӎ�,5kB%��*0�t�+/?�@~>��F�eSצ>��N��r���Xt�B���*f�{��!o�����5޵�ج�� ^���H�1z\ �Yh�[��d�6�qd����o3%'��a|�<ݖ�Uw�Z��Z
1�j7t�����o�(�[��e  I�c�r�D�"}��~���('�}��D=y#����+�gz�:P��*J�U~E�DtZ\�	��j«2��Y��kke��,�2�O��).�%駆_������l��ĥ����2��ĥŖ$ǡ���#�b��-u�io|m׋�����	���T��&�b�rL崠�`x$:�����R��'��֫���Q�i�6��1Ѿ�m�/1/����Xx�Y*���8\�^@YUc��"�����m����s�� ��8hFBl#0{�8	/PÙF0,���w����U����q;��sW�MJ���d	�Z�t�b�Mu`�FM�i�[���b|A�.RV���h�Os���/隍����>
g�-0H�f�py�I}itɝ�79c��A��ѓ�J};�ވ���+,���Z{���/�g���at�һ�!gJ7�_xQ�J�� �д^���PU�DvV�g=�\">0���o�`Eչ{?1bs2ց.��
��es�%/��t,�T��2�[)�zT�ƔDF�{������b>��������2�8ڜG#Ϫ���!7���s�������C�R�)H�w[��`E�~��U�2q�M
_zD�۫"l]d��|��!n��6EJ���S�� 
�_�q�ao�1�|b%8�;���g��*c�P7)��:�i��iƚ�#
��' �%?j��{Y�e]�gh��/}�F�4��U�Y�[�jY$B:�k#�F>�pJ�/"���+ ��̦K����ad��c_���(��Ok��B퉖<lG�8��"�{Ji�x���Z��rNB���k�����e|>��"��ĩ�F\��r���\+�_
qj~�ܚH�}JT*�x�ʹSN�(Ӥ
67�E��T
5��a\VZ��®܈��xp��	�{�����K����v^�����o�q�:ޜ�L�6Cy�W��iȺB��n?�:<�
��\X�:�><J�PF-��H[L���á�5�å��gӜ�c8��%�	lD!�YU	z}a\{L8V����!D@)���@�A���r�
H���uC�R���3F���6du�4���b����d����i@����]X$�b%b�����9~��%�f���j�����u&z��jo�S�_n>����� K��C-t�.���~���m�&��bZ��1�j�$Ŋ���l��iw��[�Ua�m�	�9?E�d���?�Xv����<,�&2]�b�3\�,'X
�����?]�<�fú��(j1�Sg��jS���IC��^�Ң?-�.V텐�� V�5=b���ԏDAD�w�Юy���옿M�8�P��cGY�9o~TѶ*��aZ�	8'$G�o�ȹ!��Q�̤f�&�e۠�P�V��֥�vn���^d� .1�UT���Ɉ�ܻ_D�B��Y���$]�U���<
� �=/�q7;�D�2����ʸ	��J���|L���4~8p~n��t3��I�-���g��D�-K�CF����2q�$[��z����B�
�%�Ar`A��"�)=�(\���FR�L�z�3���N0c��OF�۩��F%GY�(-�A�eλv8�Q��Q�Z�>ڷ��B��h!vLϗ�%���Y�I�x�s�gB��[�$��h�fW��QE8��N7Bڐ�7ֺO� ,ڡj�~�a�`ݠ>�q~��зI��š������J��S2����A��V�(!�`d�*�@\v=�Y���@���mjq�V�� �^ތ `�o��5?k&Eq�ܒ�Z������������c$!bĖ��1����(���F��Vf�`9��4�����>�x���~��	GR�.^�'5�Y퇉��Y苳]5�����e5K�/��ģ؋|_���8"��+���4�����q�ݦɛmi�s�u���3�jC?|O� Ɛ|x]״�c��f��@�y��J�ޒ�lsy�\z�j�/e
����N�70��q��d7�V6b%?\8�ɀ�i��$�����m�K�ݙ1�-;��&����R�k��Nð�j��o���A�!�_}x�B~Y2�9��>��[�;�ɂ-k���D���|5B>,�\e2ҳ�[��^��Qb��J/��9��z�w#fg�JTD@�h�_zP >;�̻*��6GT$:����ݿޓ�Q���4RX����E�l�k;ag�}Ich��?�a�/�~6��l4����NWԶ�\��C{5�����LC��Un�C�)n�sw gh#t=7A4�i-�5�">=��?QX �s���� �G4&á�?�#���$�F�N����{A��6�b�@ū��#T�N+=a����Y��P��Dg��*��MJ{��*A�qa�v��!Q��q{��E�R�h��(�����vG���1��ߟNZ�.�_R{aHzȤ@`�a��%_n�������K�9�E0+���0_Oԃ��f���Ɂi�|�V��ݿ�t��gx|��R-��ΓM����RN��8�,/�ˢe�@l[�0
oư���ld��C�3B�z��=Qo>�y�H�`*�˪����ww�܌z�Rp��B�ͮ_%��⦉�R��4o�m�U�Wp�bU?��M�>����Lp���#�=FmbP�5��%�b|����D���aKܨ�L�H��&dĿ�G$��A� n��v��`9�,	I1����c��.Y,�ʐ�8��.Xe�y���,S�u7L�z$H�M����r��ͼ(�qu)(�UF��@���[�P3'�7��
X��|�M0@ꭁ\���g��|t-X�=~3�{o�jF�*��y��3b-#��8�CiU��j>�8�B�O�3����}����h�Èb5b���&I �Ÿ�H<�oڥ��7�۟�9#�r�,k������Q����G�;'�y6�s�A
$��KeV��M�lU��� [�	M��/ltƳ�c���!U�gϨQs��\/O�X���@u�-����5o2jb��Y`��1sn�R�����S�wRF�]z�V�k�����w�'̜�����F.}�*�-I[�R4����a�+g �������8lsy/����!�n:Rmd�N^�� �\��vh���g����U�[�,̿�B~~��l�y��s��+��L
;M!�x�~��� �>�q��i{��]�r�OP�lf�)��
�b�(�ת�Ø��A���P�PSy*=���Ţ���:NE��N�@��:�� ��6G�577�閫}�S�o�>Z�o��uy�$�EB7����2T�o_�=�����
.}��y�i�}�U����y��JD����T{cfF齈*�s���=1����6������Z3AA ;���O�NHؚ�,��syz���t]�f�%��@٠���}��;�Z"���7�r��f	� �^��	� �?(�B[m�rH^���rC��݇��#6��� ���g3�՗�>1���o��^B��O0� ���O�@~r�9�/��-/��q��'�ܚ9�.���`�8z������L@_�פ^�\��l�Ɲ6/.�����T�Qg�S�&gJE[L��+�Xȇ��K��Y8���*�8�R�EP'�)�o��އ=�0X�]gb�Ȃ���YL��G�U�ۥ�&�
`���LI ��v���G�?<e0sNS�3��O�(�L$얙���3o�2?��a�	�a�:a4�����F�I�AR�52�珶����B&�p�r�L5�A�;]F��s?�Ƴ�J� ���XҲ�s��m����1����y;"���9mO)��,4`8=A⿀���s,0�ϭ����5]�痗�j�Vn*X�\��`�I�Q[�n�����([
u�&O��L��{�5�$�7�~~p?g�\��uO{l�$3�.M�W�=�D�W��%�B:���V�����b��?zI�!�k!'��,�6V�G�� �3)������jt!�-D\�q�J	�7�8�cJ��bVD)�z�%3��0��w.�+�1D{��X��/+̘���3�� ���
�m~�&2���m. �Xvp1%#H���գf05ٿ�D��!M.����?{-Oa8I�z	�׵p��U/d=�eӅ�I{#��w���9�Qj����e;�	XS��B�b���l�Έ��t��!D�	�US�V�z����X�yI���ɀ�$���+�
#T��2/��y�����|`0Hș��m
�?������U�&zP�z�'�%��r���ԇT����Ӆ�ov��U����c_
eDq.D1��UKl��<݉�xT"C!kd�~���wwQ�4�γ��jrm?$�lSux�N���Ao�����:�~���z�\kW^�4�C�� ���8��!���Bb�=�dS�1:r�	�<�j�?T�V������U����=��ґ�Rt�S�w��Jӓ���5L�poʌSQ�;y�		��UR�]��B9�U_�/;�TE6Z��~�Vks��u��b��,X�����az����>��*kB�����&�8ӗ�"��06�D�'�*���C܎��e�;\Rk<�c�rצL"�iĻ�8
V�&D��i��#צ$0	zx5��#�R�����h9��J >�xϒ��`�"8x�m���������^[E�Q��ŧPT�Abm06w[B{։�#���r��P\C���gF�#Ѩ1==�oӰ�C_�]��쿴%X��0�����@� �F$���8t�{f��+�=,��qffm��3���Յ�+du���:+��2�U���b{�� Ѹ[Nu�i�Zɸ\GW~�u��J�e�_�a(�TO�~�Uɶ;\���+Ŝ�J�_Q�G�n�w�/ވ�n�-���6�;Ma�i�C�-�4��Z{r}��u3r3;]�4�q1>�%t��Y�E���~��x 1�c�7�����uJM�ܗ��P:�@�GGR�AS�XʜQ�g��=�N��~ϻ��lTz
������`O��p��bG �u>���.�B��5Az'aU����<�a���FF��Ayz��@
G�)��ï�"Qlh �G�X5i����umI"�۳��ʛ?�%諹̯�{T�U��X}d���I�7+tހf�Mݦ��垞s7�,�n�3�H�y�:"悷�}���X��R�YU�:�`��X��5��L3���8� ���}m�ᕭ�u�d��̌|d��MѺ@W5�IƵ�ǃ}���(��{��8��jW!��f��(QLQ%�hת� �%� �\�Y�=��~Q�B�_'�\�{��*W��P��P��J��2ޗ�JG�5����"���z;k}��jG�x�$̆5��\�	��M����	*�?����T_�ؠU��[��YR	&�8���(�ΩPv��4�&n�$-p����ܻ�� ���lw�)�L�C�?kQ��6�S٪Ƌ���?z�L�� ����p������D:�$�,[�9SQ:R�lk�0�=E{{z�}���/v��H�۽��_�[hA�����D
�of0��^L_�a�JH�������f�֜��O�U���ݪ���j�sx�ةS;��xǉ�&9+̸W.�!���D��VN��Y~��/8H�n��;��UЃ��&��N7��{�#�^OD�J{�j�쇕1r�y�-L�G���GH��)0���f$�2F�����q K6Я]��;���>c����I7N���A������ɠ�����O�s�.Y A
���?�w��d�����-��1�r{�t�'�ڵ	z`���s��e=����@����r���X�0r&zS�M�ٚ؄�����������4H�^�T�TK�p�c�+�·��u��a�<F�Y��x�0��.]�C�^<o�l2�L�*�!��.��W������H-�H�Wy������?��v�Į&�]�50#����v�k�-�Z[N�la�.��z(�OH�A�<�T�"�&s�zl��dh13dI����t��/�H�4�l�}G�K}1�k,%��~�וeP�� �鱥���'do˽a4*Ȅs���WߌM��$�"p���{�}Jq�پ�xV�e.c���]E l����k4ܥh�t�|�����٧�3ד�v�����|�+�k�0W1E�Wl#��K�'�7la!Uc�{rU�}�Gh���|2sc:Hc��
a�����.u��J�׺��g8�;Uaj8�z��&I)�~x��`[�]2�}�D��(Gm�:8��F>��h&�-ϴ��I?���/j�F읐I��Y��0�aH*_�L�]�)6d5X��Le�9�4u=�"k�'��UPK���+Q!��zpY���v�^�.�ۙ���0�k@�zg���5�9e;3W���f�C�Y8�<��BJ��Wߞ�#R�Bp��T�J�~K�z��%�o��2X��Og����Z�?��G��_�Q�0z���zF�!��$��z��$�_�d?�T���A���pz��h�X�*�F��G��������$�aIco�0���=@\�����Q����֭��fk-��XC�X���c�@���v���F?^0��j���^̓(��c��x�o��M~����|�[u�k��:[A~U�s1Q����6ߗ�4[$̂��%d.��+ol�:�����5��lzN$����.�+nM����4���f*�N�bƯ5~cQAG����'ʥ�|N{�zT�.g����jW�;�ƛ��D���nCr�����H�Z�"�̅��IQT���p���bR5<��<���{4�p�<������jDA���7/��{��Ph�P6^��Ϣ�gҬ:�/�t:T�a�����&�d���5?{�Ou{#�f�0$��8|"�X�	�B;�>7N*bp���.��<ګ�D8,�!T���
ҕ�9i��}"�0yz���Q �����k�׵0�:�-��6���M{�X70.>�8��m1#h?nfp����oI��&V��M�Y�a��U��e�}^�C���-���-��X��)�}P/ں�t�j�\��݃ssf����)�ASϹk���xlm��?���	Z�ܡ�e"��s�i�[�j�V)k�z���LH�cfBםp�1(�)�r���1/��cb�K��*�re�n��M����#3q�h�`�/���:L��Į�a )�a��=�'U���Դ_z��Kt��`Vĭ�>Uo�D��@ł�m��s�,�a�ۥaK+�4�!��ؑ�z������<���-L"����ii��#��:"�|����ͻ�����=���4��Y��E��;�?L ����9#���4괊Q<{��e
��dB�U��(j%�Za��m+�)��6'M�F�f���T�m��&1���N����7�z������;�P(R'+py�����V��Y�0�sC����=�n��S)�(�&a6 *=R���%��M�S������:m���3��@�Kv�A]G6��YeE<{[넆X�
8���� �]HA'���;ۚ�M��Ư�+g��ݏ��	��M��-,�3�����\T2֤�D8�i�Jw`�5
e c�s|�e�T��Rm�} R��;��R���,A�sL�THU_�#��a�+a��XT�� ����X&�{����x�)�h�ꙏSq!�Pex$2`y�;��J	�i�
��[U�8-?+�9�!>�9�r���!���Z�հ<�MQ>#o|y���5��Ǣ֗�h"�B4�ԓ��t( ^E�#Q�}����]��t��l�D����EQ�L�'[��F<u�vX�hw}l�H�P"���\���2��*z)n��1%hM�=�� � b�OJ57;����Ը�R�.��p:k��4�&xin��537z��8��4C�FN�����`݋��'�Zpn_�tׇEe��%5{M��]A�_PV��i��@g0�v�������bpY���jܓxb�rB�n}[�7�Q�Rx;z���݊G��l�����}���vY�Q?��Jq���w{��Iaea�R�@~|�d5��/�~��z��3�J�U<{AZ ��P�-���P�%;���:EP��tZm�hAX*���ߌ/��I�; !�esUi�� ��׻qau���\|�k�u�z������/[�]�޽VA���q(_�*�ȿ
M�'DYS�;�woߨ�m�Am*���kY��n�K��e�sf 3jD�Z��1i�vHiE{ ͈��3~�ԧ!�����,D������#��lV�5_E⣚I��4��y�F�Nc����E��]���4���G<�<��q��㲘�j� �L�������l�mF�k����ˏ��(3A%뿐W�9e0[�/�6���t~S��U!����/��X�
�$ܢ��׫����8���u��$M�����X4�W��I[������$��9Y{�·>:���<��*I��t�ݠ5ЇOu���:���s��X�T|�6���;�*;��N���A��@�h���㚌��W=�0��z9�>���0���ު��=��AO͘"����Y��&T_7a�c�A$6���J�ْ5�UMnC]W�{�ܺ�734�`:ŀ�#�7pb	�RO���g̒�8��7{s��s�-5E,~�ü0 Ov,ť�K�#]����!�E"��L���`@�cU�}�2�3�J� ]`Das�8�l�{1�Bq�����ޟ�}jq�ew��\q
`Főx��zn�[Q��]db�}�y��Q�T����pI{=��?(hL^O��KfEZ��֑q@�ChH��՗I����=Q\/X�s@���0���,�[�8��ǑE r�t�B��z�)#���F��ݤB��"�̮�BV2q��Pr�r}9w:+�;$I���|��ɯ�Qc��w"�+�Դe���-�K��� �,U����	���lO��:�t(�{:Ey���~L/��S8�!B퟊���{�^ČVJ�n�%IG	!�5���lKa���o�8��s�&7ڵ1"�p�F�|�M���J��c~ܖz�t�K@�qƈ��`�Q������g��4�n��$o�7��T����uqp݁�0�qڳ�y 7����N��� �L����0��1� �9�*����eG�������CtH��F�k=�C�dC7���GbZU�v/{W�H���_��l�^�c��B��f^7S��~s�O��jv��*qR����L=��g��z&#W�K
��ED��T,�[AbPZo<i�e����3�`��2	)��untl��)���1GQ!��-�h��D�^���/U�j	~��0�@��+�j�ҝ���4㯰�����J��uI)�C�� HS�]����2^=�DJ�a�
M)�B[D�9)>��Κ� ��'
��.HR��� ��fY�)�'	������>Ǡg����%CD�b���ل��;�]cM��X����XG� ��O��pdP���y��a��Et���̙23�%�\ߖ{Kg(���S5=0��b��i{
]���q�8��@&�/��<�">�	�%d/�v�T��Ӕ7�,+g&���C.��Ld�BJ�l��We?0z{+Z����K{ҾY�m�t2����SG:gD4�یNC'ʸ��rQ���YҲ)���'?�҇8L+U�-��8���v���o���om#>].N� (�;�ʕh2���u�ﻮ\6,̅/,6�`S@1���r��f>ܪ�XΏ�jo��'��<!a�B�o�-��	o��f��΅l�z������y�O�e��/M��c��B��i��g���� ��H�M��T);�ُZ]Mۣ�e�#����DD>��lX#m��G̚�|�ډ�%_�
�;��a��;-C�?�~��a�������[S�a?�$T{�j��t�ޗ�g��W����` -��셔�iD}��!�|�<p�=�)�7���&Q����@��^8
���Q�rv�J��W�P��}�"̟K�:jE�q�(�o����8�/*��˿S�;PT��K�EB��˺���=J\��?a6���Mc���	�L��'H�T�%��R��z��0XrN��8�] U0�y�A�=�G�����E�U��u����pr�P���ύ�n���H�GޜM�n�X2�g`J(q���4�c�o*����[�@�T��2e沰+��:N�qXb�����h
�:�_ÆۓDa�+����w*�dg�46���>.q�n-���"�cWNE���s�K|�B���$�*�߸Xtؖ\�E$O��]��t�k�;��˳l@ 3����LO�1�'��k��}�ɏ�96�I%f�t@M�50/����r$�{1eh<�� r�&4��<�Ic�L!l�I�]�j]�K�������2w�bL�:���g5#cb��z��j�L����Ƨ�o�4�c�����*��"�n�T��8ߋ tp��" T�90��F?�3 �6Q&��z�F��_�B)}"�2���f\��b#�@����6�!�T�z�dvc��i����������D��A �[j��no����/ua��T�T@$�s��~�ֳ=>+�~>i��>jl���W(�U��ɿ���z$jD���ȢtT� ȗ�F
ܰݡ� �h]q���u��]<o�w`���S��s�s@so/�������i�E�$�龽�j��L��8��F����&�;Y�|����Ԥ��Cһ��"S-o�8X	~���y\��"�6���f�O�+<���-5F�¼Rp^����J�LƼ�I�����c�LQxh�wD.��^��̮�ќ7��{.��`�.�6C���fBR$N�f��m��̌���'w�����{�o�^�M�24�'L��m�i�k������ɱf�$���#�-�^C��F65�N��GZ|��6}X�O*�;��n�r���CuU�1'���9L�j�j����4�~wt�/A�0|�t�+�u�P�s'��:Ķ�����j�C�e	@��,��	�ڀ��bT OvQ-�	A�R� Lq^k/"��]�G������Ul��>���ǭ	Ԏ�z������V�VR%oVc^uC)���.o{��z�^�VA��ǣA���[��t���-!c?���B��9t�UP�oi.��+��v4WBH���� ���!���C�*VWI��24z�Z��t��Ǐ�ق:$�l7Q3A!���!��%�@7y���j�X|�$*�S��L;�8")��;'���ڢ�P�jV�5��]c�F��q0��g�QW_�J�R�eO޹**����ՠ�v���5c�y�N�[���T�AT O�����ܚ5g%��,Up�|�y<�JI��k��a�5�Z���,�
�Dg�8p3��K>��x��WS�S�[�:��?��M�48v��>ď�Ύ׏��1@��{$���[�Eg��yR�댛�(W�9�����u��k$��#ʷ����V̹Jj"�hm@���ǠW�kj���x"n���s�8��ܜ{~����A�Fω�\�"���5�?1��&�6��A2�8]�Sc�	�9Ӿ�`g�����#6��G=���잟J���ᑣ9s��M4|B:�[�1_��q)b5]O0M�73)�id��)"�]�QZO��<~��Dn7bSn�^o���'n�S8M���%�r��ۡ�t�V��$�P�#��2�QV	SUD@����v����M1�j�8�k���uh��D`~-�-׏�q0�m��	�(�s��LUJ:�d`F�ǥKB�X�M�zߒ	Sy7�#�;�l�$9�"-b�^��K2Ԑ��Y�������b�|8���{I���&�B�"��;��Dph"�AX��\�t�TH`7�n�������l��0���9+[{[K'YZ�1d:"=��Y�k�I�t0։N~�:G��s��R&�Tĸ�#�-�c�?iC�s��"Y�a��np2������>�;�X�H�mJ��c�B�:���Fs�٦�A�/~i�n/�{�{��[�вN���j%���v�!��#uDa)�
o22^�Ľd�v��F�.Ԍ'ڄ �:V���k *L���VBd]�Ibc�R��r�>]a�l�@o�Q�{`E��* Lx���`���v��	��鳊:�:���&��"_��^��$�IJ`2��G®'���E���_-��a0���e|��U�¦�:���L��*w�4�t'�:R����P��r>���s3�Jv�~�~z��ݗ}� $I�[�z�%�v��e��#�]V2���O�0]a��v��O� "�\�ZŸ]�����g-��vx�4W	!4/�UG gP)l���]�P#�	�^�y�n,�'ٰ��[|��=:��)/��vu�D�f~l��q�c��p�WT^ ��������a-��m��k���ђ/x(yϞQ�_�,4����k�dC��Q;�R)<xO����VoB.u��j�q�T?��	\�E��r�Ǘ�#�������*`�����2T��OȓQ13<�3J���D �WoCMN��~�\�V8<av�y:�����5�J&��?^��9���C��^q!�F��T)��|����C���*XI�;�R��>,Z?+� �8�M!tuz��N��9k��ޫ3�
T��+V�4ն�?Բe�f���
���Ǜ�ފ��
�@�S,�?]1[ە~�Պ|е��;�%l����!�-��",i��K���̄-�����qUpI{�8���tODt
�f�����'���3R��]OSoS���b(�8��gG9ڟj<A@��gT�(ͩ�`�ڬ?�8��W	�2���$�`�Gv1�n�
YV/(v!�n�]�k�|��F���!��(C�;�~V�i~�a�����)W/�v(�%l����r^R����+BW:.k�n9C�1��K&_a�O�:S<���O�#�e��S�"vB�2�!�N�,k��{����?�0:|g-�X��=G�&>�eO�X>>�}� �KQŗ ������]�Ix��m��6%V��}�`9z���0��|:��}ŉ&-����m_(\���{�q�%v���u� 
��etˢ�T:X�K�Qh�q����K?�@@:w�ճ����� �m�mN� q��M�����Ѳ�R�}R�'�*�\��?��#���]!��)�WN�,!���8+^Eຸf،�aCY�w��~+�I7�����*�ȭ�=s�/Ϯ�����P �7Y�g�[�l��fij���U$���qÛ�C��ೋn�b/ �t�9A��3����W��/B!t���8��t�'0-�\1��N�T���Dxс*9,�S֥�=�aհz\%I�X��H�G9@��I"�S���R�eG�g$)T��>ٜZ�I����Ѝ��+F�pe����w[����(7Χ��E������2 +3VCΕ�T���7�j�XF�^�Y�h�j��8[nn;1�6��&|i�>�= μ�2��i�D�s�Z8��w:��q�
(C1�q��s�^�����	�;E�p��y̎3ޚ��%��<�\+����z���HD%�PG5�X&,U�5X��'�$�~�Q't����*C{��(��c�7ų��&�B��	A�W�1�/�7�Z���a8I"�@��.�h��_����":���JWf�;$��B/q��I�>��R�*ބ0�.T$�%0���*��#ݡ�U�m��
����
u�@��.^k���2E�x��}���,��Fφ����2����'U�.t�&��y4���2h7��l����	ܪb�mf��Q�|)Ԣ��VcY�e�91^Y����^�gc�BW��Myu�g)z�g �>r`������9�[�<�����=�c���k�U�[�#00<vl�������G����PT��7:g��w�%�- ��Gψ��.&��cũ>���o%v�%f����|�&d���@f������� Wr�<��]��K������ʩ��
�c�bV#�َq��M��)�f���3�Ϻ![0
6ɵB|Ǣw)����k���3�s���J��v,�/S��dʍ�p5�1PGX�A��aa�G��dgT �C'9��f��QM�W���m�&����?<Ȇ��IV �v�T���h}�cu�p�I6S���2`���)��Bx�d��+a��ju3O�5:�iZ'�f]$��}37$��ã)_��1!u@
�U���=��.�%Ϙ����/�Yg�S�{ � -}���b8~��X��F<|�Y�a2k^�OU]��<�kb�ܾ��4+�r��D؎J0Z��{L�N8H��%�\��mà�^�ݿ�0e��s�?�R�]��-j��͖qM�D��7���
�&L�@���ɭ�F��\!ǳ�Fw9�~,y�^,z�F� '�n���>QX��2��a��k�U�3Wwy�
`m�
�b��;pό�������瑬y��hic���?�T����-������bO��&Cw��j�~����@���f[z�T��'H�����E
7\I3A[�.�³-x��jB0�U��)ċ@Tb�)ga�}�[@ʵ��hG���=���g$��h���g=����\Ǭ"Ѩ��>���Y#����E��w�+���[�	?+���J�Y*�c��2�H(X��C���2K��p�ݲ�Sc�?5!ۀL��#x�"n���]0�I�8�=⚔�g�|��|�w��+O=�T�� �s�`�
aH(�۠K��+���s��Q�\7�5�p�p��67_�\t�Z�C��求Mp�sJҘ��q�]�G�a)YyG���� ��Lp4"�D5�{ ���}�U���I�����3������8V�5�d�'4�!�+�lO�йt��#eO4F����*��F�����+�{ˡ����\�r�Y\��*��R���>��9�b(������]��$����\#�	_6J�G���_?~�Om}�#'����������IT˥� �x	�塣.ʤA��y�Ͻ z��G`�6W<c"^~��Q���ŷ���-��k�%�|��XZ�R�u��n0lX��r�vm�X��- �o�W�H��>�o�Au
���J"��M�:������� �DA��c�
∎�l�Y���ͻ�۰c/�1�y�+�K�zO���GX�e�����p��o��Ђ���NR�Br�:vћ�;]��wk�1㎲��L�Dd���myՌ(O����hl��7a��6�����ұC�g�m����]`�G�٧ou� �Ab~س���}b3�!>��E�y���,�I���!�V���xPMޑ�7BƽgOh\n�H��\�Ć%��D@P�X�K09Un	��S��L��571D%�4s��m���W12��㌂%ej�"3K[�'c��K�+EC�?@`P��Τۚy��嵋��̞����L{����iN5���Mc���_6��J	�\b78؝X(3���ߕP��?8tK�p��U�E�U�N��1�{��f9%���=���:o��pkO�\j�ϕ�Љ�(|��˺�����R`�mn��?���W�>�~��K�JԷk��1�!�{<�&��( �qC�:�7e�"�t�|��!�l�`S����̳3�:�s��:�}��l9��z��z������-���t����N���Va�^�'����"Wa�@$C;�!���
 2b:7h �X�v���%L��3.r�V�r)NlIخ��}�8!�U
�Z'�ۏH���pG�Mo�X���j��׿��FOmh�?��rl�*�yx �Yb&��S@N֡*!پ���R�cZx ���S��%�<=R/��3�������7��v�4�Y���n?����T�-���u��U�F��(`���D�@�E����lơ�n��I� �ҟ/a_UB���;�Z�0���s���x��[S==�[�)�.�J�*�W��ryr�'ˈ�����	�e���`s��e2f���o=�|�{9eJ�:I������JCyN��ŗ�d�x�U�y�#ϻ�f[��41�]au�*ـ���s�~��������d��^�M����|0�MC��'?N����h��� j��9��K�1�ǫ����� �Ƶ.t�7c��\y����I->q��_����Ƹ��f؀����VR��n+`B��_pV��R�q��+�u����|���)�L���c�O���p�
\M��2ǌ��uC�~;�E�̖~z]�ۈ����F|R���(݆����!ʹ=2��XP�T��W�.���d�I�n�?��%�
D���XO�a��ua����Q=3f���mGR����S��d�B�� �T�l�V� Pb͠�eb��M�<�!��j���*bO���Ao�Ho}TLfR�"��ns�J�7T�I>�Z�Zn!L��n�����TU�d֝z��_8����T����B��/O������?�yqh�o��fs�&������$�W\^�7�$.6H'�l��.���]�J���/S�rSd�QA�@v�U��L]�H���a �GW�:���>G�)`A]
m�5Y�2�����	2Z��y�D�M0��QX�����g\+���C/����r�hO�^��ɼe���Y��3c�K7rR���j��ۧ��@,4R �w� ��]�IU~��32&��o���t�tD��Մ����.Ώ��(Y�_$Bi��O\rOz�@�,�T���ֶt��8�[[�pai�@��K�8D�I��nyY^Eƙ6;렑u ���_w ��)�فZ_v$��
h^p2*�	�?��JMW��������>���x��qjs�\��+�����o\pϸ�M���!0�зN�bB�};�#".A�W���W�� I��w�ۂc��i�؟���]�ke&�'�@ux�C��p]�9���j��J!q8�����K�Q:P��Pg���!�j������g���Owh����|���C�'����0(��`ݐc�!��7h#��dשDOk2���.��q*�Ji���d��3SE{~��u���H-�r�e�V+nR����iU��2�j�Ԉ�͞#�6{-5�G89�,��0u �Tԇ�"��v̅�Jk�g�C�V�+=��V�vFD���E�y��yu#� N�lO��W�K^����H0�~r�S�^eW�mK5q��(*c��]&tZ��4$��q��;�~�Mr'���g��������==D�\̸��AR&Q�B�U�a����Vdn3�e1]tP�Q��!�l��wg��9��W#�<g������T�Ry-�j?d��
z�5$���P��M�S�2,���2�k	���K����Y��:�Hb�L��Fh���* �6�����߂�q'�d��~��Z� ���%l�K�TuxW�)'��輞�=�r�#�x32ȗ���zx��K��]�����;mnbj,t�.t%*݊N'�.�1��^U7$�g���L�����4b��L���a��͞�3�I/�q�$~I���Gq����A�Ӱ�l���H���̢�VQ b��lQ����lUđ�'���aVIC�J��7��b�zz�n�0u�T>g�va�x�ǿ���*vp��ɻ�?�
���4:���Lh7����f@7K:,�[�y�l� 3`E	q�}׸�1�� ;��EJ�z���ye���mk%]�k��[}�C��ÈBw&=�|�j�cܴ9I���9�E��Nq��,	ԪO(~���]c�A�Za�8h�a�^�5D'd{0ħ@�K=�i�@#��֑��RP}q��tx��m��e�&i�E$ ����D~�߻�]T]c22��>�e��G��"5'o�K��	�x^�z>̋U�Vs�_%���,Hu�y [,�#�7s�+H>��2dG�B�����Xb�9�^w�i�d��A���'�|����U �n�b&�?S����̲��Kof�<р �K�y�R��(p\��uB�1� ��Sb��1n�:����E�ߙ�H�|��Ț����|�nq������+}&��u����M]LXk������� $qv�͡o�-��f$ٜL��A��?��e��׹gk9 MmZ	[M�C�=�2 ���؀t���@T��Sc�\�jE�ɓ��艹 d�G�%�T��-*t�����C`h<P$�q������5s�RG��=�RƤjI��Ɲ	�7�z���Qg�E�[����/!�N;@���*[p�n�04z;��Cl��;`�p�µd���z?@c�$x�����j9��'�3=�|�Zk��r����҆����ԆD��G?�iUr?�_Y���=�u?o	]ӂ�0�6(ϧ� m60��,��P���=Y��I��O7������^�Ҧ%&�����3p�u��>	CL��/xF�0�_��'�����Y�n@z��x!�oqX0��9ݦ���`�{/�bEا��0e���~�W�I�XU�<�Y�"֞�K t���*n_"�^$��%ajY`fBM�@�ң�z�Q��Bf�� ��6k���CI׻R�4�H߀9C1�+w<t͈జ-ֿ/� �4l�p��,H1��x$�m�����+�g�:z �l}?
��°�5ȳ4��OЀѯ�Є퀛Y���#� ��A����/�v5��c�}�oS9s�8���{�C��m�'�����~-����$�I^Š�vM12*v�㜋�V9��X�C7���n���=��q��Sz�OLl�Vv�dV7������L�X�Ke@X�R>x�*N��ȉ��$�� ɂN��G�`g���x�R^�&���}��m�����E��[H�\'	ἡ-�:�F�϶��A�,@�5&�F�h���7�Yk�4��~�����n>��F�*=�X�.��N���A�$�4
�D-�F�� c��,��=6�𦲛�刹P�*S�Y����g�1ϭ$a/�<-aY-�-�k-�FOY��T��@j�`���pg�K�3�q}�8\�m��7��-��y;Ol���i�{��t]v0���ܰ���2f�W'��K��T�?�I'��.O�q��?�O�]J����
N�E	�K�"D�/���{A>~#%�/A�[j�$������K@��'+|0�e~����^�P�Pĺ�g�������P9mkB����qå�m+�Wgy�h�0�2<\!�
*i(�O:�F�*��J���s�&��k:+��퐨H�j��;2��(@œ��$���p��rJp���������T;X�\�#����4(<Z6M%���ir��j��a��s���So��$���h\WCS%{%9�EG/ n�����}%�L��s	Rm*D.Q�t����_tZ���<z���k�7{G�ҩ��K[���E ��H4��
�<�o�%�Kn\���,��!O4��,��
�JH�I��	��I��iP�;c�߃�/��V���W>m5Y�	!�*�h�|zz�*�1Y+���o����������Yk�"����u�x��r�W���'�a�A��qz}�b��8��Gy�[7���h�V���ص�J"�)$�(74�o�<�.��~P�9'(��i�'���'[v�lq�����������3�eI�&��k�k؍^��(uL�=!�纞X���~f&=����K��5a�r�+P�9��~2��2�f�I�@��EhPF�Lco�?L
����J��h�,E���~�0�%���%I��)*P�p�ɉ&���2_�h�9C�C����_GR��*]E̫W7�6d�M�rީ��O��H���CZ�e�hSâ@$�~h�6�3f��#Q��ű,2�;�T d��,��Ω�4�7��x�������S �636��/С\�����^{�.G�� z�wyH�.�8�!^�,����qX�.t�R�R�0/_v|�!���Jѕg|�sT��QͶj�ߐo~0'��p����
�_g��28�UǕ���J�0Gu_�?q1Y�4?���U�A��c��\�B�==�+&�1��W�p���Îw_n��?��Jd��9԰�������k{]4�	rH�CB ����+;/����}U�pE耛j�?�����yʐ�vTX����t2�_����	Z׹�x&��� ��f��V�Z.\�V
�U�s��X��1v2��uc���_����+�{���EP�$B�Z�lċx��;��m,��Bd��M����*�E�s�=1��J�^B`�&�`�(��O���s�"�E��zC�A�O��NR6����Y,ZEdշ=�[6���{�x�����@����	���7>�^G6�%��6A��ݮ%�|��(oqE���9%_�T�BB3U?�gy����=���|ܝWG5��+��ݛ��7(h�'\�=ZA��������ݷ<ƿ*pl��38�ǉ�:�=G�1�5�@B�*�%[�O�����D/�\��H	'.�R6�bU'����$60�����Z�\�@c`F7�{����Je����+�,e�D�F��
�jx�|Q���r/(����wƦ�$�(�5��E�@>H���{>��2Y��s�������[�kRs,
��4�Ñ���p)�~̣�&�i}���gd6�Qߦ7�f);��vy:����Wk����Ʒ�d����x���)cL!`�,$��DL>ׇt1�og��H׏�e���?�����"d��0�p���!�t��[`k��v�����������ɻ�ڐ�a�)v�7@�u����WN��P��}�'�L41[��� Pi�=��T�B^ɇ
��"��n�����mTy!5^G
�_���'����d�y�z�LT4t��q��f)�9O)�!ґ�B����X��t�����k�Q#���7˹����o�ק�&Z��S��e��t��?��"���2l�Aw*��2��	̶���u���k�d�P�z,�9{No�z�o�ߛ_�o��jܽ�;�c�pV�4]Nom{�V��W�U�� �N���̱5�/<��d�%�2_�$����H�\0��K �����;N�s��Ax)���e��k4�?gx�<9��%���^�[k�kjp�@���c*��GՓ����m���Ъ��-0U�� �T�P�vf��F�Z�,�����q,߬��o:�9��9��O[%!�����ؕ!�`�j��<���kQ�F��x�����0�U��W��߂�aaO�i�%�-,I��j`G�K�l_n�����O�Yjn���Tj0ޑ��G<U۶��sOj&G���\i5SyJS�(�������N�Ȏ�A�#5˖�7~�4���l����(��rUWS�A{l��=/��+7Mk�@E�$���ytdW��m����.��hop.��)�!�Ѝ�V�����b���A��W��pv�sw�'
��?��H6A!U�Ό~j��K΋�v�\�������gK����ڬaH7�g��(����:���R�=�*q0��V��R�h �������|��Y�{�F �y'2�5��A����mI����l-��`��Q��&V��e���Uc��6<op�N`ȳz�f"R��
��~��Գe�Tf�?���ZG��:I�΃����6Bwa��qL}W"0���|Z*k�s-�(����g�31���y��dӡ3�
��p�=�ҠL��O®\6Ko�]��[��J�"����������������5������1�9Zr��.�4;����g�����pK�ˎT�+P�z�\����z`�n�m:��8�(h�jf��X�:Uxk�}�YD�����u��o wR�,��de���[�+�.��n2iex��<�,�g8��Q�"Zy2����9hۑ��Z�7'	��9In+��uڪq#�r���2ZD�D�������5_U��S2��aO� $�8���mw-�m�|r�#�����9#�D���^F����K����y,�D���T2s	
ײ��0O��v?
-���ta���c�<:jT�h��G�!��m�
T�*�K��ҕI��m���!S��wr���]BN*��L�Ҷ��7y�[���fg����I�QiA?�	�>ʌiX��ϕe����Lt?��`v��Dy5�����e�Lr*Y5��{UlW1����F�n��RJ��eۣa��F�
k4^�pK��	 ��2m�@��yB+P3V����k/7Nӱ@vg�]a��9��H����2�ri����k����3%� �Y�����g׶�2�t��18�����oa��<�m�Q��)�pX�Ck�N���4?)�9�
ܖJ��tM="$�����bt����ąEݑ�������=-l�D�\Q�&v����>�����d�x���Wu�.�����5'��ѳ�����.�s�79P.�����J���Kg[4hG��-�����t���(-)�m,I���'G�d� Z�2�7��X})��5"7��I��+xR�)���[� ����"�,7-��3��tp�U����Fsc�����'� "���kT{�pg$1�fK-��]�U�y&�vo2� ~\��I/Y�l��U��+���@S15�.ǫ6_�>�Ȟ�8UD r������W_r>��y�}�OM5�t���0^����YIR]�=~5��V�7<yɢj[��;	�LD�� ��ڀ� 8���b�9mO�Ro�;�V�n�˰[�{;�bc�.c��n���ء�M��!jJv0������(S�Va�H�LH�O��h��]��
����So$���^ ���V`d H~�`��#@��<��gN��9�掊��v���H��g��w���@��[����D�7�B&\�
_�ј�XN��Xс	�ny�������^��g`YT�t��$X�+�I�`r�%����y1}^�C%�=�����0��2�E�BbR�F9�e�J�0�v_t��Bҟ6!sm��9%P3���Y��A�p^��2,��x�����\E�+�em�4�N[Ĵi�#��y�O�R~�@k�F��1�rpv��1�C5w���6Yr_*$���jD6��J����Z��>�������^��<�&��4��]ek���hE��(�a7��:���t�p�f]�A�}ٟl�dhs��qѵ�S@P��6�!�CS��3^`�
�j�ԩ�AZN���l��*j�&!������� Vx�*�
]�U3���)��ղCȿ�EZ���	qiP:�w���+�{K��$��M5���-2w�6+*��L�I������P�������kΘ�Ă�y;�`���I�O]וc`A��l���u�c�e��a0"��oV!�q���s�0��p�����/����~}�u��#�")�GCI	`L��y���<��e��]'T�4�����l�`�B���t�E�6��ђbub�A�@{
ʸ��/���(|�4�ն�}����;y�k����Á� ͥ��7j���([���(�\c<�	<;� zw�&�R��
Õ�����ϖ~�SJ�,�3ÿ��jei�ar��C4���Ai;`�\�gfɩҎ�:����w�osZ���o�z�O�<~cQ�&Y��V΁m����	z�Jf_�%�^���uY��f��<3�*6&콚��) �h/����T~=Dw)_L������Q���AGo��|ѯ��]�J6(A�m\�9�>�&8W7����)\��G]5V�L�k�/I��I�i���KRx|T7����=��$zރr���û@/sT��B�=s�\
L{�ņ�pk�m�?�`S�~�Ϭ��	�DY3k�@�'����2�m�S�a��ƽ��9k�k�Dg�ϏN��5뭭�d�ݡ��pC��6�^��_pY�{yB�n���gd�]�#I:��KQ�S��Ɔ�n\�e]��2��d�?X���#5bT;��\�8��!�sS-�/��nRm�I��-K/���{�C��̽�������@�~����8T��&��@��Ӷ��������imM�i]ۛoʺm@c�Ij�P��f����ܻ��.��e��-�=�	�����@d꯱�tQ������]����F��*";���y�F�AG֐3,�cG<�+�8C?H��q~m�kޞ��-�U��{��2o"C�s���C�g*�~:cyĂ�@vY�����T����UG��
mB�S�ٗ�Ҫ���}����(�x����:ԍ$X3HUC	c�����|C��r�Ǣ� �j_.��#�_`�_�>�e�I�0]�]~<+P�����U��P���F<?���.��9�Fn�P�.h�Z0΁��S{���P��蝧b�qWP��ADe�&�{,y%��߾&uqe2Q�c�*!�)<��Y5�MՏ>�&���ȐeK�L���,cY�$�[0�A�3w��x&�{�J�s��+Z������2B�J��o|�"y{�����s�,â���
�G��+.�[���vJ��qI���l��1i.��9��X#�ԇ]GZg�+��1�i|�}�m�1 ��"/٫?N�R��J����!�����\�Z�]����.r�T� 7��rŕ���!Tq@� Ʉd�HF5*�FJ�붩���Ë́3ls�݄J����.����p�f��d,�-��y;�޿��1��l����[��W*�e}|��(=f�����V�D�޴���,�;)��?*��*\ɭo5y�a�c�l�]�+{�A�%��J�ƈ�:BI�{��T��c�\���:� ��g�h����#�4��(׻\Ͽ�̇\��x�8�o 0*:R��T[]��t�W�tv�]��#��>}��K&f�a9���YZ}[�j�����s�Õ�٨��3n%�T}Y�W5j���8X�W��:��5�Z�Hs�!�!.�	��V]�b=�����)b�T�t�=MT�H�E�<95�~�;A��*(9�r ���5��n՗i�؋z�^?�߅n�j�f��(�#�_�|�ak���O̽5��I����H%��0�T��uPc|���|����_��|E&9|U�����e5ST��7�wϦ�`�|�|(��٢6��+�'e�j�����A�N\�?�7���Nl�W���
�U� �}mK�KO+�'�;������p�-ꓚt%B���*���te�*mY8�{�v��zO�� ]�s����hf��@j�t��t�$�O������|�L\ �����	�����й ��t-ų���j^��e^�,~P���a�>�,�%z��z�؊�_���feA�/��Lj�$I[L+�[q�����n�<�u��!��vZ@�B J-���_Y�\y�oi��^��k���d���<E6
�3?&�I:����c9�G�"�o�����eT�Q�j��s�a�i�ޠ-���H�_k�A�UJ��{W����K�p��*V�>����2��`�w3o���X�]��A��)���t�͙��_��U��4_�]�}���4��.y�)���I�
m�Np��NV�x@���b6��0�͟�FS4�̡�}8����4���z�jp�J,��W󫺙�[�����;���i����H���Lx �� �d�e,�xm���V#L.�y�}�ՊB�0j9�8ٷ��8����5>8����j�]]��d��bB��	,=J�����~��"��?�޸D��}5�;Y]����#}qn��q�Wע�>.��;gSc��5�Z���zl����
GWdA�a ���w���iɼ��~+�Ո�鲳r��٘Y(�̕v��N� R��(HY
�Y3�iO}��z��Y
��ҬB��%���Z�5����Ǉ�M¿^����Y����M]�{��:)N���Xdj�/�S{��Ϋ6/9aq�|��]����g�{
�4ծ��A��޲���	��ۦ��������\f4Z���F\7u��C�4��b�q�j�.����	s�;e�$�ɏ����׈3� �
��Ŕ Y)j���b�Zͥ��f���X.���=B��$�49^��.U����o�݄|��5��)�Ǆ�D> e�)w5�/��d�gp�j���kY�ͅ��O7Oc�+�2��AQ�#@��d�"P�_�+X��Mϋ��dҼD�Hk�}�׷��ʋ^��\��!�ڔ�*��Ȯ��e�D�]�x|�����M��p0�6�C�9ٓ�J��!�?E��A�C�w�!��� �$�?1o��_\Xٶ;�up�=V�Թv�wwa
���S-G�/��s��:5���44�9,3�] ���`�僆j��>!Yoɉm��k1�{��0ϕ��/��\Q�F362��1#����딬`�=ۼW&�I�/깩��/u\j�vF��H�>�3�����$r�p_�#(���
�j��W��@�)A��+*�U��6	��e�W�'��i�0#A3�0«���3��F	 x�#47�ꕡٞ�H�i���l�����t[����5��N����s��WكO�^,���O��O�	7��#!��MΏV�0z<|I�oE6\���-[��WW-�m�����7��
maV�X܄��/��s���Bx�3~c��pc2$�rfa��%��c]�Y2r��D��$�o�Je��8ӕ�T)��C���?r�c�Ч��ʴ7#�2�<gR�+Q�)���F�{�f������P���뼲�F�e��I��Z�([$�0���!�Vm!�Z.��_�=aW��(�8v?k�A���Hlؔ���jԦ��r�j�ù%nAz:2	C9���F;0���3�v�̘$]�2�*v<!��%H�L;Z�Yu�=�bO���U9z�s�V�łK%`�M�&� &u�h!���Md
��Nf����%"�k�W�x�����4ƞ)�1%�܎�1�]�=&U�4ɇd,���cՁaz�G�e�z��ޝ�W��<O -�H� ����J'�{@�c���܊���(��&px��9h�|���C��#˓趇ȴ�z�K�e_<�2��)S,ٷwx����4ߍ��!��=���*_�-���@1�P�~�}�7� �T�6��,��	i�5r�K��L	�l7Y���m�ij���~��'`��@1���V.ȧ�m����u$}.�E�晴�u0/ǹ��@�t��u��6u�L���`�1���&�a���(���G������j'�2������6��a^�v��k����x�#X��H��Q����d�t&D���\����ʟSO��]��`�_~U�.�F�R	3
%���!g!��*
�}ő��6�L�j�݂(�a\���S�x���-�Ia]!D��g�ҕ;��ǶPz����)�r��`��g\��ǇAL�$�i/��\)lZ$�jo�Of�*Qa�z��O�A�
�%����¦��3*d���*�EP�c[�l���]�<uo��$�N��<-�U5n�!n	��eʽ����_V��<��Я����=z�GZ�Y\�91Nd��{L�%�y7��c5�4�.�e؟W�2��Z�x�2�AN�O������l��6�Z| ������P��$�/n�$A��xMM��Ml5�rp1Uz��U�v�,r<C���=���Z���E�D��d���4?�c�[|�?����2��S�l�c���ys�%���z3phxXqx�K�s��Hǒ�,�B���$��eKj�fV1�%	-��h��2BJ��t#0���1vgJd�]�Ń8�;F�6�YiH<Өl^"f6�g6�D)<s���u�iu�5+A��h[ bDκw��z�#L����3xG±M�8 N08Mo�t��Z��h���w�x��!X^���+���Y��I
y�)�S~��D�W�#�UQ���mxaw� ���T���Cy��߸=D8���:��Mˇ4��o9l�K`�v�-���Te��:H��>8�>XH r,z߄�=*5��=\V�����8,v�k��ͮ��J|.��<�ءMi���j�R{���v;r0U��_��u=���Tů!ﮘ!��Xf�e��Q��s7h���{�Hn� K��QD�)��x�� _0���E�!5���,�W)�4��I���gެ���V�����v:p"�:� �`b�/S�R�910D��i�������n�#[)�-�h�Z�����'����GhY�����Z�zm~�G���v�=������G�d�4�x����`�Ŏ�!���G%9˸m��ic�~Q�1ȋ�o*�bnmk�qT�׸궈S�
��<;��.e�X�����z�,���[p�a4�����d��>W��-����wSRy��&A���'1�c/fi���sV$�n6��
�E��O�B�`�$y��{#�����=h�X(M���)����0lo�y�'�>�<"�@(�����mN|َ@�]]:X'ؓ�1�r*VvUM7|���/�����R��?�U�&B���Gp�ݟ%J8C��x��V�h�_��hP {X��3/�U2%�1R�O4��$Q�����T�����g�5>ĺg،��0���������J�T��~�_I	��G�JF�P�n��Q��/sQ����d��!��,�J+K�u3f��^�7W4m$�{��V9\���G������P0���B��������N��к"�c����l@��CK]�������t�aܚ�kϋ5
�a���u>Um���]�W1pd[b�z�Fen�A2���LQ���,���D��k5��naVc ���Coy`��s���gy��]�t|��V@�J;��g!Oi���V�3�9Kx��1��-�\���s�uM�I�<��l��O��r����v�C��&���t�*j�Z��It���¤���O�.A�7v��9[X��(7uP���mi-���_�����.��ZBeJ\D��E��[����7�w$���F ׯM1����k���DDy�*{�K��1K�]r��X��}/���q�I�B9�+�*=�#	���μ�Bp�U����U;���������GM ���m�z�h��he�~�b*n����+I�؜��$	�o�9�eul�wW@F4�ܳ��-�V���M�i02��8c��q�2ë�æN���=^���УoIZzͶ*��(n�
���/��c�����<b�Ș �:%M��0T�m7�ҽ�d���@��t-�D�A^Hu��%�2;>5�+�����8kQ;�ӄ��5da�n�p�Y8nq!i�p���#gO���ho��;����f�~�RQ�YZ~���^�b���8�/c�v�����Ц���[�5�����%j�+&\%d�2��u҅e3���,�ԇ�d����ZѻKY�A�yb&d.�4�N����.�/L��O�K�:�1���f�&J><���*ێ'A��B���ݓ.�}6��N[p��6_̴�B��[�.��u������p1 
01���dV&���t塱؟yA��L1'��Bu��#X�z�;k2D���N�_� �^��fQ̌ǥv�P�.�p|D��E����!��6����3w+h���?�N��UT:��$ +S� m>��ҡ�g��ӯ�q~�c���&l��8᱈��������"��&�o�����'�B���:�*|Ow��iw%k�IJ3:j����Uu�h����RIE�:>�z�����!�¨��x=+�U3;KW��׶�����$���Ҙx�=��K��"���r~�c<e=T��r�TQ.�	' <u�Kf��t�&U���!�=.x-:
7�� �h*��ѿ����n7eV4��^������>��L�W���к�ݮń~:�cL^&�HkT��7P�.���!�߰��Y�Y"���
�6�k�0q�N�F�%-m�v'�S�O���i][�"{q�O�r��q�H��a�
��:	n+�RƓ��d*��`��uHJ����\����sh�q�4�"�`��ó��
�KV����	��￤�B�Ҝ
�5����2~���/�=�O�Z�<�����G�s�I��]��|�y,F�Rx��V���z] �ݙ���@���NT���p� Z�ю���_���=��m��7������\Q���X�&.�{7�4Ul�ixǱ�M[#��&���{[�*�9��ڰ}E�|y�{1�0F�<�Gf�R*c�n��C�+�!�:dA��y��Dd��~���^�[zzrv�x�R�����o�⑭�ZT�*0��޹`�	�Y��Z���.���9#ҏ7��-+�>����΋�<P�j��JX�<
��&	(�~�E���ObR}kf�����V%�]#(�W��Bƚ��IĦ����?�g���K~M�c�d�m'>�@��+��i�ʼ��Po�f	���FTJ@�ۨ��̤m|���M�Z �ڵ���������@b��j��
L�EZoE4l8`jp@_g��^��t3Yx����W�i�v�U� o�D��Ҋ*;f��n] ���b/���7^�,�C�B�^�D_�MR��R���@�u=���>����ۊN�G�i�2�S���V�����=�h�)f�� _"�Cr$�k_�����d�}�.�5F���|k�<R��n�ͣ)��y�0�-~ /휹t�-C1c� ,���Y��J	���t��J�I ڻ�6�j��m]i����v�U��,�����bPw�
��|>f\�AM!vĚ�8��qa���M,W(P��ա1i����/]�t��v��KQ\~6�-����A;�ts�C�{��>5�Q�c�ﲼ*��d�O6 1 �lm�I&��g��3M���i�BU[��T� ������%����Qw@Խ��1;M��ra�x7��K�Ы�dN$ S����i篞xJ� h�ݲ��`�ܪ@�~iF�FS V�3��3<
���G�Bҷ�PpJ>8�?,PK�Z�?�	�(��@3����"�F;�mjT)$S�7�{�7Z�H��3� �G�
���x�u\�S]���/�7]�0�"?ڮx ���UFDzP�T$�נ�T%7p���:O���Rm�Z���Q�&�?Uzq�GJT�⫦&�(�'�`�'�%�:#�f�B䜄6������>�Tǰ���59U*��[uU!-��W���6#�>V�a؄8���s�i(�����i	�HUI����mz$*��7����E����?��9����`̣�m�Z��Փ���vn�.S���Y~�Y��R�QL֧~���&� ��L��� �JB�]�؃�6N��9`�$�UN�n
�'��}��x3��M��^�~�z��N1�1��z����$HGë]�=:ӷbP�:����g�sIvE����E�~���M�ة�1�`xW�M�1�~��J4��#�����2Vn� F�WB}?�����ݙ���B�J�×��]�B"ɨ���~��B왔��pgM���5��b�(�}?�2"!	�:Ig:[�@C�{匜��-l6���j��ZK?|����rO��g��S��_�CY�^�0�B��-7{�5@��T��G�@��p��� �	2203�5���
7�+e�@�d8�\���e,�?-�I�쥪��GM�8�nm�^��݄I����`KZxYj������`���V�ņ������5�e����YMe��y�J�L
�����v#�v�)0�Z�#i�Є�l������3u�z�hs�z��� َL��Cv�Ɋ4�7<��>��A`g����|J��$:���7��:
����� �.��^�L���Ǳ�/Y�9l�nJ�<�2��e^ۯZ3�����o��7R�zu%�f�h�#pC����'[=�غh��]b�O���r CE��%Ji���9�`Z�>d�U�G�L��Oc����L1ʉ��D8�&�
�.�n�(b� ��TŒ���� ��z�7p�MQV#���S�f��Ґ�Y �%�ޱ��m��Y�L�(�VG�m���KA��g��A��!�ӭ�xߙ8q���Ú2�v:�3�'�M㨦��xM����rai�O
*����hf��g��!ώ�p��&paqyT*AA�,V�*z^,��"�]%�JO��;Z�?Q-`�h��E�Q��\f?��vnV �!���)J{pAw `Kw�~e� ۄ�cȅ@���s��U��6i�P?6���K*E�L��-3Ƣ�GR���ز����
9����j�� mw��Fѭ����Y�ùV�/�K�edL��I&"������!��t�����N�P*m#��>��eBr$�8���;�������a� �u����nڠo��Y�o��W�0\�������ɧ(�xsڱ!B�8��V��e����%�8�^�R,��b̗~�j��3Z� ���%�/9�y�ed��q&�Z������P�:8,���W�|S��������y�)o�Fup�%���c��޵q=�f��.�&;�>c;:q^#1��Zu�<ɸ�l�s�������n�Q�-��9~�S�n=v�6�}���qϧߥ��#x�7����*�rv��7z�_g�78hP�R�(T\�ԞWD�şNd��l���|FT�x��~N�Q��{����rT��@o�����O�����_qF�l�$��KFg�X�po�����7�7�M:����2Y�����i�Ihi��sa]��T��1�Bቴ��:oL�q����!b�X�X���K�è�MD�ة�^�7�"���ސIb�ifz����ρ?;�T�M[�4c��K�?�:�)��j��P[��ޭz�qZ�1���^�Cj��5����Ʈ�X��?˾��9��d�Vљ����OL�/_l��,T��Q�b1�J�MW^�>�>`���i/��w����m�0���X$�������A��U�g��^�O�������̇���U����ՎT���}@B��M�M
Ƈnt��T!��{Xq���?��:#��Gn�cX �y�ꋷ4�G�Ot4�w��b���u�wؕ�AU'bvb�fJ���HE빷��W�? �g�!(r��;�mF�������׸յ�V��xǐV���?��U�A9��&U��>8��^a�x&���y
����ѝ�5E>y�A��)Al�n�������O`���J�`�(.p�����@��j%���rΉ7j��b�s��k��,�������2w�K����|�h�@�Źa�f�B��NR� BT�����D�K�!�/c�ژ�T�/7s�>h�b���f������ꠕ:RLUט<	�����t3�_l��6;{�T�UɻU,
�Y����,�Nc`j�(�(�H���3����#��j�5�dz/��tܵK�ԙ&� Е�d>V���K'�2�[�̍��-�mCt�1�B��@�U�ϛ�b���Y_&c�
uK��i+�1����$b��#W�L�\S���~�7�1Sen��`l�k๗e6�Uk���S�20S�U���#������m�t�Ϗ�)w,;��Z�4ň��SW�8��q��R �K`� ��ݥ�*4}������Ǻ��9e��	���P�)�]�(������d�^�6��;Ϩv1b<�@�*O�S���N�?�6l���rxk�tLr��V��&"<Q���M�0�0��$��U�:T���3�����~!9�]4C������<��S�璅��8�C5h�`�ج̕y�S6`�c�oB��-�0�V@dE�q��O��H��,FGYQi��{B�(bSm����L�A��]���Z���{;Ħ��F��l��j�o�ć%���W�ڨ��It��7�A�dn��>V�wOy>XU�kv#he>�D]	�d`{�{���{� {T�� �p4�MjڬZ��<��^���tl�7�];�O�9Z��p��� �n�u�>�yA7j��k�jx!�X܀Ք���A��#�w�<_2~��q��ZJkz�IG!�B���H:����?�7��29_G���G���!h=��(�]{��J8��M�۱�>�O�^z����=�с��T=�J�rCK�I�K��uzMg���^)v&N��2?}��a��hxZ��F����sG�5L7���D9*hb��$�$9xf��`;&Wb���CN�.<w|��V)��%!�6q�Oh^�v�T3�=�w&=�b�P��p
H8Ԁ,�y�t氫��9G�����4I�bb�u�	s` ���}yo�l�y7�n�(r�m@�|GC��k�&���Ohآ��n��OB���p�U�.���fp��M�+-�t�
�ICAJ��j	#e��VBK���O�VM��DX׍,)�z'�-?^<�ld��(���-����<��xy�Ҝ�â�B��bjq^��P��
vK;!�P�,�wJ��q=�������|	�\��]���s}��T��J����<�T��I��k���a��]z3��t��"ܛd�a󲧣&����M��:U�S�B '��=ܱ�]K%��$I/vLt	n�Ψ3݆�D�L��o���`�=� ��zq�Ê$-���@�3yY�����S�R��n���=<ɇ��'t�&�2���G�^F�[(�N�6x��	�6V���0*sm�aQ�x�?���d����52:�v}SI���K�15�s�*h�i��9��Dk=&������p��`��>�{הMc!5]�������
��A�}2�q]�|�k���0�-2X�2�@�E㻃Z��O�\����P�F�C��w^S{��-�c�v�[r*���őW����|����f�0�� -�w���aܹ�֯Q��
m�͍<s0k9�M3��lc�����(��FC�s�Z�$�& @߄��CcX7o��~��P@*����{��gvD��R��	'7�ϼ���/-���]�?	��x.
�N�m�$�Ap#� ԓ�?��(�g���Ж��d#�_J�$e	w�>�oCZj�!�U����D��<Η1KK����C��6E�h[It���'��r��^6�Ž�g����V�l١�������5��T������k��P����YqHg��i�4�=�z����4� ���FM��=]�0��ҷ�u[�@�u�N ��<�g������1�U����Ϙ&��D�pa��&��V��?S��(3m`N1�t�v��[R�,4���E���~���#�Q�Ǭ����/9:@N8��n|ũ��:ތ׻����(մ< ���!d�-�m������<%�g�M��K��+�	K� J�S�X�\i��vCu9+�i8D�W�ؿ���oZ#��bʛB��w@»�gm��p2U�z�j��oiK�8)�c�t���5é$c� �(d�i�O� ����tSB�b���e��s��߿6zw_�ܯA�W���j��5�J����b���HVn��V���r�
����Qҳ�&�P09�����p�^�V�a��|9$�v&̣�uI	;�p����Q���2뫤
���+���'���&��g�ԎG�G�X�o��;�w���&6�[�r�S�K�x���F���*�P4y�K�� ��Ωb	��	EL7��LtEby@���؀����{��ۤt`_�[$!�|,�������
l|�8L����x���n��4-8���[og�9��I~9��g����{�	 0�Ҧ^@o�V�������l�t"���H��s_�3=6���)v&���k�//�P����ġ��E�<�K�%� ���s�9��PO���f3�P������0��:�FqA��`��� �f��h��ƠavFm˶^���_��&�4��K�z��=�RU.�l&{>Co�d;��p��M�p��^lڅ�~���1qsW�8xT�Fm��V���.!�:Ĝ3cݧw��C�^�q�=Q\�Rd�g�e�,��Rק�q��qO �K���=ഛX�$�xf?�����WJ�|0;�F�&��΂�pusoPA�٪�PCM�^s�$~�"��sM�/c��ܗ܈&a�b��E͹aJ@" ��f��:��L�,"�W5f��$��s� d����u)�e�2S��	z��#�c��<-��1��Ɇh�"ד%��8�_���'�F;E=3��e9�Da�"��(z��aF.-���K�Uv��U�Fj��!�w��Ӛu����ʨc3�lh�X���ă���&f�o�m����N}�6��M�h��T�����̹��b�-����P�ڒ��Z"l���B���4#P�����X��qy4���n[��t�����Le0#|2�?����.Y���.�@�N�G��m�&�ԷDvW���E;��TkUjRFB9 �)/�w�����%}�5�p&�֦kȍR=}~���m~�s1��e- b�����4�܀��܀o�l��Shw*�Q�oiHf���a��S_ٲ}N83�ڛ\�{��B�[z�HE�[^M)R5-��nY`����-dF*ĂӒ� ��6~�*'W{5LA����L��!�[��[����:ͩ�O;"��)����a%r�--��9�/Ӊ� ��Ju=-f�D(�t��3Ҟ�0����9(��`�S=?Zh`L^�n�짙-$ͯ;v+ۺ���y��Ygц�dѫ�H�����&�}�'SFˠ��a-�@�B��f���L�t'�ָr|g,��^��x|�^{9�խ �6��g�ݗ|�c�<*4�Q$y*�u�I�Fm�dSJ�h�`��L�H^��c��L�SoT�α��?�@��
���c�Yqv���),>+�}�~�= *�,.�v��)O��o��4�SWFu��M�<�k(���[[9:�<����>��Y�z�U;����}�t�� p��棄������II.t����٭θY��rR)�b�:�6�x'��L�D��OD
�E��S�ΒqBף�,=��������:��ų�w:#���}V�0�-n_��ڤ��/��{4�h8^)t����:� �$�+���HMW�R}6���O��>e�V����u��;��1`t!$y��_���f�'j^]����-y��@���t맲��iڵt�6R[���k��&)w/J9�S��x�[$2\����Z����|9x��ǧb�ׄ����-g�S�ETG��-��uYl���"/sr�'��[c�uɚ��v�v�t@/��%?-�g���j{�nd]�4T��k���!]}KG���GVˣ"�Aoh1�Cy�Ç��q�SI&џH���k��|��1
�Jl=�U����c���7S�gjȹg�{)�b�Ԗ7c�1Puy���������{�;8���P��bd���B#�l�6sU�]l=���rp�	���q�9X��6�z0=���������YW��0�^�~V���p-���[^���t��؅��n�<}��<{N����F�ac.�Fҷ�-F�j�G�R�;S�p����2�Qڷ�S�����0%WW�5a�?.x�p�UV�Z�l3Td�*���.����+л�?98�E��u����ߗ~
qP3��tt��*��s��U�&=�����y!DX�� �3����=zjY)����e��hd��x�?'�����G�=���*-v�0�- ?����^iK9��7$�����N�� #����Ґ�q�@3Or��'�X�(��=?��jj�I�'��ܼիy�v��������v�, +��m����hV-��7F��^;�����X�p��&�i$�	������hR3_I��VS��,����b�LB���j	u�˘�[�UH Ug�7�C�|D���p�y���xNT�e%�y���9��~�`�j7����	ȹR��|�řF����p�?bg[��GhK.�w{Go�\G���h�b�cE9����$�9<}5�]��j����e8��������IqqO"r��z(�y^~i�S�C'(v�n.[G�$y��T"�=Y�#��X����0G�UwZ���փ�n�Eˮ�tX2�*ژ!+�S���80(g������_�D`��?Lk�LҼҕ���Nl\�LȪ�zt��WU(��x�-��=BQ�I;�ۏ=�~}��sg�ܵ*]ZSő��Q`P��҄��� �l����'�/=��0�gd��,ş9Aj����V�4�g�dv�K���W/c[����zc�3��L���%�S��,Q�R�(�1�1~"�d�(m4e�{h9��\xέ�
�I���jك������ٚ,�c}�m8��{.�����T��Y:1d� =�Pyw��k��Z�PJ�CZ�w��r�l����͏j2;���Pr-vU���Ͼh&������9y�B*�WI5ח��8�8����s{r��}�`+��p�u� v�|��h*M�pZ�:)@n�]Y7^wɘ�g��Ӧ$�'��dW��o��ۀ��2�p�M���	M��h̚bP�y���ޏw�)������. �_F��T���\�Dy�FI��o����>�aok��d��9��c��
ZG��4�j?�>��NL��3��/.,p�{�l�Ģ�����!f���w�W  �LEyIP��V������{1��ԗ�:��^��K	�����Qq�n������)4*��<�s��;'����H ��["�7�=a��|8*�<�{�Qu��GG��Ϭ�OsX�M8󞘚!�=&���'C���%W�� D�Y[j�]H���"�/Gݹ���?�詴�G��c�2)Tq��j�5,��bLK�	f�1_�.UX[�z�(�o��C����s�{b�*�r��5m��%+�<�/*��E��Z��&��m�)�S�J�A
�e�`�b�柮�ݫ�ڜ���;X�h���Z��?���7:B5.�z�!w�a��&k�h�/��A" g��Ł��3H���/���U��3`Go"x�<�0Z��GK0��K؄���a`�_�s(*�@�'Y0;��1�Ϧ%����=��Q���Hn�eHV�D����FK�a��?2뇻}���<范�Ġ=Cm}ۇI�I����\z\s׵���R����=��C�Sx;L��g�h.� {{�X���/��_��|��f�X~�ƾg@yYLf\�I��#��xPv=͗݇_�#B��kߺ��ԑs`I�ml�Ƈf���J̈�ˎWo��(sY�Ǟf<��J�6�&_"��{����	��a"��9���M%��ݕX���GNT96F�p\i�����'bE�
��|ј�F%�Ҡ#�i�0)�t��F<����m�!r$v웝|�d�>-6��E��:�"C�cF�^�v&�%��ʑ�s�	zrxA@~�9T�&@�f׵=��:�<�4?���ᢴ�B�|�S<��9{_�׳�L�\�Y�["_E��;N��I����x8tN*�@=,�M�	���.h���.�9��g����=ؚ�P�w��@5KZT��R>MR�fϫ_T�>�5�����˰�>�]�{�1vK�A�]v��^�B,�iu�ޖځǍ�[a/��k��`�hʨc�[몟�9VaЮ$5y��mn��r��s&E�`.1h�#��O\d"+ �&���m��:�~J~�R���ۛ3�����G�>Z��E��ŵ��%������$�\���RwTu����6���\\H2G��{�8s�Ӕ�OF��f�@e�:��cS� ���.�����N���:���ב�uM)9L���9^���*5/��>'tsF�3jD�]���H�-���x=0*�q`���@ׇ�4��
�'X���p8M���L7tыiW���Ĥ�d��lC�����������3X�����7x+�5�]��p���~M�
�|�1��w���©�.Jw��E^ӗ8,Xi�g�ꯍ͕$3�)P�.�b���;z	�7ޯ�,"� �{GFk��T�`_ �����1�)�M�����d2�r���ﳳ�f�]iGث,����Tl[��0$wƬ^r�wL~
��꫘!�Q������'� k�Y��#d��f�r�d�-�!1��Q�i&�E�<J��D�t~2�~��s��O>�gl���s�]Eċ'myn!��7��b�����Zez�4����Uw8��kT)����̽P�'J���c�!0И�)*��P`|޵`w�>bq\�'[��;
IԨʲ{����xi����IA�'��K��G�J��y_�y�RV���� :��2\��$e��{���"m����T��t���]2U����Knா�ᖛ:�f��!�w�qN؝'tm|�)�s��P�#f�����	N���A�@���sݾ�o&A���*�cj����� ѝ�(X_K|hu����ػ�Dv��^ӯ���)�U0��Q���9�%2fG�Ɔ�#����gf7Vn�k� Ԅs)���F�z	xC��Ʌ��f#e�BXDb�u�K�����X�ࡘm�)N��!��,l�I���0�N�� pVCm�I�O9�?��-]R*��)d��x �S��������r�D{��W�޿�Pۜ�v����^�E��v��S�Rz:]�2��R+��I}@q�;�|uu8��X�`�ҡC4;�!��``͘�x�2��及$�-0���j;3'+A�ŌcRs�@�9V��V�N�݁�G�v'�;��hs=���Yg5_А�����0� ���AFq�H�SIÌ��>� �^�Ӵ��R�C�ڜ���{�,B�QE���g�f���lݷ�H��$�.n.f���Jd�z���m�QG��z�c�
u�i����^�~����o�GF�aO֍^�����w7��YCL*ЧG`!z	$�\��j�Ѿ��=,��7V��esޓԤ�Nŭ�Jp��:�C����D�?�f�,��b���׸D��{���~��0:&Zy5�.�'�����Re��uM�"�|z�Ok��0k��|�X�،�7?�%6���������g���Q4�J�������~t�LbĽ�i��h��O<M�.
r��v�l���4�XN�HS��ls؃�c�.�뉏	㌠�����:��B���5m��gS#�u����+ڞB����,jN�U�4��9Yf����8F`d�w���^Qr�{wݧC��0(������B`��~����1SP��0B����M��]�������qw���r1� fD�mk�Z���T��G[�Y���8�Nt���:�ݣ�>`�9���Е%C*�4���.�L��gz'��d0ΡIQu���l9;���L�k��˱�X]�_�N�D
�^��UN�����*����C�3�)Ƚ�4%%���4�� E#��YWY��]���/bQ��c��~�X ���\�$\5�/����,,c���R�bJ8��.�hwtkJk��v��+҉�3�^�M�=�:�t_��pk0��EO�a�e��w�y}c�F8Q��d�F٦���9&�~D��v#���w�ŀ���Q#����h>�/D7�d��������c.���x���pi�R��a�f
e8*#V�{7��x�$���a���9��>e�*ت��j��Uǽ��) ���̟x;��.�ع�y"E)�A��ˌz�.�|��?��Ψ.�B��%����t��.�.�)�D���ˠzL���9k��0��#BN-F��^s�����'�l�"y�ݱ@_G�Bqw�K�,��BzN��XEvݺp-j�[���i�eF���#�E���'�'~�dl��e�j!DRa�q�~`�N]�,M���(��nr2́�����D�gB��l���v$,��!3r�j�Аn��Z�(R�����<h���õ�<�k�6pΤ8��vV�Սi��k��I��D�Қ�s�撲��uܬ���T� �i�Nҽ�����݂�)"�q)���#���´%k�� 2k��߭2h��iE:}�L��f*y#��֑j��w<��5���Ã��~Wr�b��|(�/S�׉ ��ka�g�1�ͳA�������c��n�[�8J^lj�6��e��k������>��<���AU�~_�nH�4�[P������f���F�#�.eD���.��n���@�X�k9������r 
�n��[���}I�*�l���]����<�)��t�{(���Q:�/�oa��p��,����<V��YAӶ`*�Ӛ8k�L^�
X�ML嫨W��� ��ά��J(�eB��}�����-g���E�d�48=�3 }2��;C)