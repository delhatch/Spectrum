-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Z1Iww6Ie9r+56r7a4zZa2nz2Vqi7rl3kkRCTGVOgfFsVf8Wpl3UZ6AJVwSW/hIb06KCUBSkwe2Qi
FCdrWuaPkp/D3BPwzB8gf9IIwIiw8p8rX9Cr0SFEo8/54MZkJyTzSmYTeDtQT4bwbi301FJrGY8E
YVJSEUAoRhmaPdlMLYw7J7UeukeN83Vmnp6trdo4lrUPVoxxthLdr14Ewe4V2l5LWAaCdSaksfS4
k+ZwBgz5IFeqPKUKlQmVxAveVFaxK4LIwx2iLl+Zo62tiCc/htxuiD8nWgqV4s6dKi30krm4tl/T
Tauib9AtHJN8WUBATRMsNEbEqjNJj1q6PiWoMg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
iw05Zos8mtNY9RG+ozF7s0dJ54lZc6ADgfoEGgvixKyd65z4WxuzglK+ZK4xDSMpTYhQ5XHt/6Il
4MxHbDb7BWM4GKYv1G82MKv4x6vQ7+hOjiouOCjJndspqW/7quZ9+BFts3ADOXsy9btQzFOq4qhP
CdXTVrBejAWR/FXGO8KzTmrL9FvnT2PSr/pOm9cDhzrKcZdb/MPxXe7NQ1WypmYkYJ5D3ROWJf73
AGiSYWzd6j3xzfssxPljOoFvfk9bbwuJC75/wQoB8t4dcpJvEAsfUderN8xhTibHDsEdfkphjgHb
7U+0sFoMdezo4ziDKz2zux8GfPNQOXjTbgwYkXjeK9s2cnnNDJwkcU7QMnRZFNSKo7FPEZ9o3U9C
CBXj0U63r9WE+FFE5DbrWr2uaz6qMbZwV1yYUA0PXCzZWt77tRBYhm56xFbz0dOsiG++Qvd7M3MX
C/bwUVuNRc4ai/mK7MKNLT0gA8FZHwohN4fa+rhNP+FYxJ6UhkeQO4Xd/fcaOOyNizcZ1uZl2q2/
L4sbUIUKqcs70vp9tGSmNEl7EjCBheoaLMNbsFrPC9JqRVxcJ0Z6vGG+rdUOteSxeQPDmJGObZE/
BVqmqEaiLcTjsTvX4L6dfgiJ6Gk8RL4xpMyHzu/4jVPIk0bCpYEB/owhwTtJrrJmLVNhAsxwU5BK
cMAslJkZufz+lZElx6WuLrvkKaTyyKPyocgDLFReiHxV1c8NOVJ4pKYzF3Gd7+H/E55/ZbULNmND
8ZyPAW6qCIU33nmy3UXsd4UcAr5ReSJtfSJ5jUbpLX+2uVoEwQnjvYUSXegl1iQ6uH1ffP1MsIl/
9OLh/A5OHZcBCoyan6YU+JZbYvzM+qsT08AVsv6pP9LvJeg57IVwUBU6SwmwwmzPZLBCj7dGA8bK
Oo7L7sCU+t8bcPRF1CUDRkXdoRG5n/2JojoDFuUxlJBGi6amaZmOSv3j/iPL9ztCgE/szkc+Aexy
sl4kDWvnOspIsZGAJRk2eBr3X7eQ8dS+Gc6c5u/s5FagBY0J4zND3ciy/uIlOU8gycmlgoHoCmRv
u0UPA90lucXPt/L2ukoTRlI/lgmV/hJ+GV+wUyj1VGj4G+UMZ0M6/eARcsHOAMrTwBEu5GHUb0oq
VcX+gJBOS42l/g0TVyesftRg3v2fYqCoAZoXsZpzYvHFR3CK6bpnYD5LgKNzIJ3M6//RZPENVD7f
xECzFrO55X3IRsjV0StgCzN88QfJqQwhRSTK8ZLJxxe78WdwJQX1SQKR26ZFk7S4lR0gRVqglIo3
Gw92itvElboIDFI3l7QgEcAgLSh5Uf3XNBo6Yi3Wox59tOzH31dUgMI8DMCIK7oLEa1MoKmjAhn+
nMxzzgmpuIAeSYtuwcJdwBR4WUch0xZENOFmvZgR7E+0MUWSlf5a57OdL+hJ24eNPSmKvZo8lULE
QMXAAO2QVHjpoPUQpUL92nV1LZs4tMnVW+Z2oh+J/OHo1c3CqUYb/L5RV+jZLPxOH3J2R7zNLnuw
JsbZFNvHWvLe44Bucosr26T6TnChZaanLknEQT2u6LcLQN2SV90mYgW6eyjqF0siWlhqcRPFWK1V
FHbmUj9Q/O9jenV8siYjMBj/zfly1Rb3OLj1r9oPuViVxJCh7NnWWGzTr5FtLvahnFFrzh0vO6vk
R1Q/AE3HYaMO6Vx2auREob4NDO0TUh8iXbOUUpl004X/6aTs93tQ0wstowahICd0pzxUJYA1aLk8
ZAPsqqBfY5t8s365xojQ7iH071EOrMWfz8D9PMdtWV5OQo7PTEcDoGo7Wx+/No/Y7yVux6P7J3i2
5k+Sa5eC5+Pytm2SMnj8MHangkp+66V7sAFOEbsNzOxwoe0eoO2hqYfHBRZpNpoK1W+iEam1V/Na
jWN7fogyRfWIKyWbdS6fSw3DvmfXUi/vYQhE1qJ6fKDpq40feGstbHJjDwgAbsVKFHNRZp4+/ZfA
2OXDtPuFQ1lt6yPyV+vBX+u0Pe7j8EzqdBs4ADdjbzq8ZhhEvTdOy7FX1E0IM8jWQCDL9rLq7LR+
773BMJ2oBEagZyoxlmHgCj1ESnDGBUy833nZYMgtO4E7QVqsnS1Pbylvou2JzVlzy7oMAauhmxV6
5yuK2nZo41uMxNiNI9ycuVOMTAgGfH+gPPAXc9HOzs+QJ4ldeKScte2gK37EXpVl8sxzZriRXbas
jyaTqsRABFHGyL1YCyD8q+6JWH0K1VuQFHjXVdSqSXmrwhq++A0HSEZHm1oXTRJXKWJZFvgkwhoe
XYU+1FNbZUYCP/bfyO12lag8
`protect end_protected
