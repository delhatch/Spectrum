-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x8r05uVMuRpGSfldmSVB6bmo+X187mYcEFlM9VC56468ffyEtkH8aTZGC0Js3tZjkVN88Cfhr4hl
5zp33OmeocLMicApd4A3UapNaPOXBb2LpUCQRC2BdAmzGe7j2Hg++LuPeEwGUub6mMXqURj/R5Z8
0Hjx6hL0vDOmydHt9xCJ+zPZq9bda3zya7PRleEb5tBr7W/TuPOgFyCFpRmXEX5b5f/g/cYxy2Ln
3sGTLamZsDpGkc8G7G/uPxzA/3faUS3UVx4ui9vd4GesMi5oqmn9aQuGTQq98KLc0ypEaNjTSoRu
naJFotImckMR+ud3endhtiQgzEh/CeD28BEYJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
GTSgwjC+a2Ujr+VVId9MxzIzTHBepczJSiQyMULfMFxxgLLWUerLv/H2oMy/hHYQAQzoyiINPeJ1
mEkSgImmR1x1jYl1h/Uu8HhSGEZGWRlEC1D6LcpiY/WEa8+Ssd8QK5abBHNWA04mBid5Lgd5uKjL
iXZegoI1XqEPWwMXBkOEC1sEBFBviKPLrV/OTf4IzZ5jS68FsVAclx5b10KUarkR0EU4fojo1EOS
mT/rUL123svXycLXSQFuWM5F39TXo5PF/ujJRrOT1P64TsUdoeqea2YNb97Wyx7M2LFIxaVgn0Ud
ZKO012FPSCvXJgur6cW6DC4yTfCkJPLpyJ3obInbreVlcLDmt9dGt9D0UjtIMRg34NPF1Ysh/jFu
WhRMRXPJrMBJXUn+PVa/inNPS1dAzQgGAbtN4bPPPMLuJWSq3PhBv4P8NXKxsuROS+oelIrBhRJN
rfoiAJcz+K5WwY/DbmNh33ieh5m5fFEZrWBXr8Yq452pB4glLCtyr0WNCvPOUMugDmhLlZInzxHQ
LOwHPCgJH/kQrox3YKElcwIPPBgFMLfTdnXkQEU4DNoSpkmRoCR1lfO3VP11wrPcO/PUCJDIS2W7
/IvrTCwkc+kvwkflTWb3ahpQ1pQ/VPHdlABglZm1qGMFXBeyc+NPAlLb+IC0+bHQy0OjXzdu5V6l
HifDLWJSw3JI6TmBlTCOxrC+53FmJ0kWWNy+P6mZta/lu9PEq0P3sZId9Jl5oaqg0lvZHwwmnXFs
wecC1PtOQVUODyreFr5CbHm4ZaCVqGbG1ZeeOi6LEmeF1Hjgms8JXdaZcsHHgpqAoN5TgFrinMmP
O+Jm2l7YjrcyIx2R+b4hfM/bPj/BpwsonzPglAs284pk6f4yuPNJVoc6VJCM3wYMTM6rE6CYDxAm
mYD6GZPORl0OBmCPXaz97AdeXzeQW/om/QETD0qakx4iQVNpbAaAtxBxITTxUbRpXQnWzt9yQIkm
msXcyG6C5hr9aK41NrG+xrEvx1frNL5I5k4bmI7VILqMTflzKmqM0kYWpj1hdN1OHhRWzKx8ox8S
j1qtW8QHKlRzeD36Tn/167bQ8MFEN3PR/QIxbfHQ6GU7oLqSa1GHm+6PMlzepu0LdIgpvNiqXFUe
HkBMnH0PDX7Ev4lviaLRNx/fTf4j4ehumyah9JpLwCFtYu3bvjzP5TQA4gn0iKqZz3iUYfu5LVlw
RVOvrgTib02nK8OopS+Cc1ioRdFEaIdmZJKmWkowcriTAIKkeH2g/gnF7AJdtxeTQ+lzCLvBKHBn
rVy3vc+q+uyh1Z3y+7+/xDpiwu/HH+4CBCFemhsaQjFC9Gcg0ocE9sATau1GMgxFCbcgTuvHET7z
BWZ0P/DKnMczeSJ+dEgTGWBilvvDP9bTuj95i2DDhUPIn4+jvAOzMT6EWQXmFtPqopN6MVY1uJpy
Ui2lrtAFZTG8RHPqCT8lv2mZvJLeljVCBdQG5UP630dNo+gDkA7H8GOADg1bgFu6WKtU7e4r2AAL
yU/Mf1etnA5vSF02HJfMUepq6/S/nSoscFF/7uUnGEVf7Dx9av8YKUZq/QpraccppA8T9y5+hIUO
EkAfaRhlJrmoH2vwJTvfiQ2dGTrLKU1wGeOXuEq8cePTO1zxxrKbjG9VtloRZrG9B5PaskM2vCqk
To4za+ZqUdW/aNWGtJ00l4+EeevLoSBFbQehXhqLz8ZzkIbXjTAiKiurNu6QIYrYiQDIGwvfUrk5
TBbLaqfk/hH91cHAJPQALQ1LTZaxKx9mxFA7h37RaE6PberPaXJLeDITFCF4ZT3XMr8p4CK33mgH
i51h5690tsN5qYJrKoMOZqdmTjV0c91hbKoMFVkdJxomIePs2BTKKcfMqu8DjYJATZmxdKDe4hkq
2M/sKYZLhrxxkkwOP0Fh0pbRkoGAG2VpfZb+pKM61qf938eM/VU5gJwj4xoaHUWYBOIVth7ThCuw
4vQWiad0VC8tsnxWIuXSqKylkKkrGNlAGwPVkCYUgIfjMIKJv6/+nY6yhV1Emg+7Uj3VsFjWdJWw
iFFov5xFaWNM3eiYHDx3yh5Qa0eitLAxrTV+PmLGzSaYGdrnQvkAB4z3JJubfYUJH36UPQ8n7nes
PGGWpNRf1auNzm52epImbgwUPbyAqpVodCt8Mgic7DqSPz58TFHAqkfBTaXKHsUTEa71ipF/XS5Z
+UnjSv0JCebku9ADAd0uIZ+II6HVMn/oyU7BX1hp67YltA8flmQnGBLTB6WlI0pO++lqlHQNxDsM
ktbsAaUkHmDGBcKKosF/B+sE8oVLAWo+poSYcEUS5Udncl2wJ9SaOB7uG+dbzSouJxy3KzU7rhhg
tE3scULZN0fu2+gvMP8moYTeRfzER5vBTPfI/qxdNkAU/YHJttN6kI2ceguhJ0hIXgIUYqDvPd+r
Bj2UN/ocm0HPAOir4Xqz37HPWLwJ5rewJsH/Mz5h2mkzu+XJnxezSZcrfIW3v8as2FasS7O83/ES
HXxPuAXbpO09EMuiWrHz07o8sHo1Mj8vBiHaATr78MjDrUzwpw014o8FUholxxTay9CH4sRkR6eW
CFR5QBfePNZYcwxamETUv4RYo7AfrXLHnXdRl1iBW9l3TA8MVtXNecLJBn9rj+2cwBzN/sUXk5PB
oVXSthO2q5b5HO/BoU+8TFwc5lKTw2pkzswzgF1L7h7RHPAhrSfPAFym2W7J6X9EzPosctC0Esdz
Khh5oGU3W+dVABADFR2KUG0PzEtrqUTY+cnH0jAe6PeprQnKuDy2t6DvcJZ1nJuTQoxjElc7EkJw
MULKlPbi5wXSTvKTKHhhEbD1jcJK+icjw7uLII1gGl2pAYLX2UHu14p+UOEz+NTO0uTQkZsL9nb2
5riynXdE/9NkoAoCwHHuzX0t1Kmz0yxAreJ33PKGZRJaU32EWR62oO6G45Bii9bULuAqR1Z9LvXl
glawUWr5JwuUfpCe7QShzXGrEKrT4UhcW/6EY0K9tBf6GxqkraFpW1g3lAv/co1SpA7tHNb8emuw
vU3DjUT7CMrwlfmeZBFvoeAZ4Y+C/oZQP59OXnSgoIiiVs1Herz1P/MR4YjSw02QddfzgCPqM6ju
fZoyvECKK/N6Drm7EA39jkMtl0x9RFGXa3QylW+0OvPC9XDyBhe1De6H1QnrsSJ3VH2524n82LoN
j+Loi6PSZqCLaXkoa1pvhU3uKtRZ9C4JQl4ZzanHRumk2vad5gjU5BuxcdtXAAnMr5A5sSeh0y39
hM2w0Y2bH3QCe2aq+p9jY5HThoujKOH118TRLATUT+3gvz4AIJj9R8DgGlkR6Osddpiu5pSVSzi7
M98V7t86gScDGxBgu9zWKQCl4HFwhLuF8GqUMJIyYTGPEtr1Y8KkVMCGDbnndT9vv3Bx+xN6V1AZ
pusRocIepp1mf+GPtbV542e55f4Gra1pYiSuKrAOCacypWAYnfTRWUl4hYLbGlFYU2HFFaGinv4e
2YF9jmHsdY+RNjaM4Ran40IxE7KTxtejKmqQlCEgmPlfTKHRMAup+lUSiNr/pcT3zOkJo/5VTBmY
hII2gFczoCSURYCA9RxjnnURFnbe8aH/eV4GYEMBa0BxM0/0W6ZPnyj87LcXS5V2TxNO4M2X765a
Wty96GuIxvUJbsJTLKMX6NNI7EemQPzOl3CXI/7Ze1Fov4Zm0d408fdKkMUxuqPkYcDEE1ig2U2c
b++bNzkgdfiJ43XExK2HddXZiY2cUABg2xIEzV5eqOM/TtlbX2UoGmyo1kwog/5/jS8XBUCmrspn
5XXVttm1dvoEV3gFq01mcTUEMivGFR0tk4cQZNL3Cig/W8I5Sl+Cs9lZ9D2675544HC4tb+Ls3dM
b9gVp1RlVgAb2F40mF2Yk752SYAgmKo12Bnypxh/CTbycy+MC48HlcWq+glxgX9Df6EQOER5pYlz
CRL6dY6dtRKNW95kBbbgMaKnBkduJQr0Jmwmnv0GnvGw6Cjbt7fevEjqP0xjX7+ngTPYYN/se2rY
aAbFd/lWtT/wrNdTuXDbzvnPleuQY8qVByD4mlDUfMa0+kcJkDFMR++e2/6/IGoTzUFr67R2mT2V
xp9+Q2dtvt0mgskwQBnH6LaNGy1EvmK7zao9/peQsCtoe1J0JtnpOgHEB/yHOXNGPUqN6Dacyukr
/N3jCR/lmhvAME9ZGeQQFBhni2fr8Pze19tt77/+afrSwnaeXR0Xz0/YbdNxSyzoCk2kwLMGfEKq
1kdEVATaQJ4pRtZnc/eX5FIf5fEaRfxZRJlz3ndHmJq8CgKdKeCA+pbIqacbV/gXsikuIKj+fZ8j
YyhGhjkuXAmVO6QaObIl/f1xSk/rbS6JA0G0cXkJO70jgrNwgxKeyRCmyEhxCuPgQjr36Mw28JXQ
IlEoPo90/p+xuLQaW92f839k5r75wTCAr8RNENEKFiht2yKGXE0gZLuZ32WuKmIUwYdtU9g7Jnvd
7BesPAarXJQythwcm/5C4zAkMYlrtZZOf5W92LXJMnrfYNPIIml48wgV8U8EkQd9XFfSAFsVJEZB
vyLtLgoPSK86Wa/b0xaXs+nSKscbpLAHdrUW775wnTjE7EjgWkg9hekKqWmhWz8uGMM8V4lM7Gqa
omJTRwEKMzuBTD5hV/eUhyD/B9GKhL4CCiWx0grQUFds8d3UL5USQ5D4wL7+CQBkSNZO8SvJZt0p
vdRthCjL1DHC8mbBwNBUyrK0WUtwITBWxdNQtos5hVzDhCYlpJZfsXk4H0W5oftS8yfYPUhvS85p
4yT2ogLOlf6uHCSlmBo7t4sIcE/8+nP0ukCXitx+7VqM92p4a55U4bEUl98y2ExIuZYqdZGiTZ54
CJyO+aVg/PD2thaiBAgtnhjlahYYxnYkEcyIVDvEHk6ZFeMxLWe9cPCp2OgUjNF/4OSE4Ot9TIbl
XFS7ZVwXMN9o8ImDlMfmIRZtDERWP/fqYIdGAdN9EGxyX160H3Msvyviz5rkPgjT2lHvrymEikv/
YtnBpg/p8T3k5SwFNXYIUa+YR4qTapoQ7nJFfJ9SSt5E+1MluIUq/rGIOiugp2JYx8fCC+Xz+O86
KCOnFyi7rVIgSdx2gKSvE1jJnEDAu0DQEegoo2T0gPAHnuW+8HEctNS2GDg8Qv1ShMaDFG2WVArq
wlfGd0Q04qLwIxPilVNzNmJBPG1188bj5pYexFy4is5tzCKywwXEDEpso1/GIK7KgciavcYQ1Xsa
oN6omc8TGuqUv/kvxMAhq+ir2Q+Ex4gMz7kGI4n1iRYiIHfDOiL9j4I0svBkzXF71aC0OrN7o0mu
J+WRH2D4R89m5rOVMueIZtAaSA/3kYFutZglsDskMeFPHnOTTIOHzQIrLqXEaRRG6/7GB0V7Vx2D
8NWu0Jn19z0Mi+jBq/fASa0IeN9QmlrBT2gsBFWmWaYn1gXOaXJDMHWhsmzs4IYTZ2ZN4nrA1gy4
68JLMHm0XaeLg6nnyMFAcUI9Js1sAzbIYsYcQtBBFJPtYxp7yAARlh2Aa+WrvUE8075yrtGeN9Kb
wZlSdULOfHHSD/buf8EnnokI3H17de+2hhVz7x8fofj5tEdO9ZjMdAvhA7ErsKj0LtNjPdeUe4kc
Jgm7FtrgIrgfmc4awkfSKBerxsbJvddV5LJJMawgOt7iOy8mcjj51dMOS66qON0yfZaE5UoMSlWq
gqLEPYyJK75RpQQxWYn59muyzBvF398CCJ2bi5m5E4lSC3DsZ1ry6KMlKuVyob7dkUMJrdi4upS0
tXZIqOrrDZ+PyB3c9RjbbLWSIl8kLQsqw9zsNhn2EH2/Q/k6VIOK/uNFtvmu428MnMTlPuoLdZLH
FNCQDl0BD26dd7N0gKXO/E7xRj30JSabOoI5CN7Ovr8ZG7o3y9dxuhCBWuEIqpwLD5Rl50xB8JKq
RYVyHK14wlHZUEy52csRohA3HaPoSz7NuhDiLN8wXslSdFuDLTNuzzo6atCKYCoPv24I7hShL7PK
sDANj8hnJ20qj84/cTX8R7QpE1NATEPWQ3VXXcpNHVzToTVdxGNbEO/m2EfrXjHHsbXD6wQuUwkd
FLhmSDOD9FAj9bnncH0CgrFGrZZ+46I9l8eEHlZv/WkZuImkxTIOYOR+v48NiqwB81eXUmUvfSEi
03rxE3AuFtwkD1ly+YYD1HoWjfFzFrXyzCxbSXfBIz3UAdNhTg2yqsLm5F14jUvfDL1S7Ne7pTWs
uIfIHNQRvvu6+LQD9U64reLsY0zIQFqHXjCptIumSzL8tPYQOmsOgFc1k+SSPoSlxSNmkW3MPSUt
IludCxHhvLEqmK4vaRnKd3PA7Nue9RVL0bSEbbx3KZSqjkB5nK4r228BKyCSzofEFLspOdXCF+0e
Uq6cXErLrHTVR9igQWWH6F6MS9OKt7A282O3O0qlzbWOCU6dAJoWVAWNbVKx24ZJ+NF2GWu+xg4Z
6XzmPVWGYJ+g0TnRM2jk3gLN7A4IYolHE6fbAawwZQK0eC4D+d4URqbkv+It+VntV6jhvjhlidMk
XJDZhwYUDgrf7i8tMQMWoGrgO8vgQRtuS1Pq0peK7BWsiDVPNwa8N8T7soUIiNVLh1eKIvPYjXWk
AIqMvyxWkFNbyYcG5Cf3hfjlW2+MVuS67k08sjbwPDjcGS4Avn1Dnerl7e2qmrelFtUHqhKTZQQu
srbZodGW9WMrUkqX4QiMg4KY+AqpCHo7N/hRYpz77ag+dikGruYtv9wnqZeSAQWmPZ9td1Qb8Bb0
ozHO4AtmykVgkOmB9d5k0desh0LwjVx5CaFn0+iAy1Ocm0fxoRzle+fv3Y/PywMJGC+NuPFe2s3G
JC2jSXFsVIeKAwSqlyWWE6J5Pd10mwOcTcgrWdvC3g3ZzAwHLMJtNZmWlS3pKIgWeCXPqT5AAd8F
gYI64n4znOc4NWOX3lPrc7XUP+dkPJ8wafElfDym/JFvI9yIME4r7tHr3mdbVD8T99wlZ2hlPK9S
Pfwc+/P7eyXYbcrAn59FqEnwX8rkEKtu9k29QqgphgAG/moM8ZLSmFlA1HJecAj48d99bnBgJgx5
Z8AiwbmY7OU2bQg67Dlhk8SEzy5DMzFEpe/NAWtSgNKG1SUCadjnIKhESX7hV9edMB1EswjMn6hu
w5jhvA5kGE4mXDK4rZRG8+Q3Z+Z6HCE7HeUNm2LuYJm8QrFLEi2vSfsHC/gSgMHpjDeZY4ljMcU6
BeCLs5vh6s8eSDbsjihKREj6Y4qsQ7U7QUqayxUtPfVKU4cQ6Te6caOW3QKogRvgniHpZvNtZD5c
1hnADNZn+6TEB4GYdCWnTqyv/rDPjgqJdK1lTPYdciFDerenvq9UA0NM8g5T1jfKl49ScmasijMp
WIWHaVTWAak4iVLsYd5i/eRL9kNOr+2JT9Ra3ufLcKzYGuYpPEfIBy/MoGpbJpaDkqCHzzPjnHiA
FB5a1Jc2UG2P6Pkux0VqfKIr0oShu6ybfEpvPPTJkVDPTP1MdvhD0yAi2Mv1ubCWoEka/FUITj7s
oDwaEea2kI+DGZU49kD9vp2ISi2sKut2WoU/UWNmtKRXTNG57HqDB+wCLtUofTqUfbRpPkCcxhdC
SNkBfZnzVhA203tp+uoUXGKaUL9aH68pYEV43GJX9A+eFUFWy+8lz9uktPv8WyBTkqaoJWMmdcp5
5Qdrn6gdjzn3XL18Bbul5hrOk7HXpJ68SaBtMarDvTF55KpN9AabCrF9CqL/8pok7R0USRFrl6JG
rco4+Qd7Wz2+KBXMKmq0hFmuDz/7Hn9Z/pjgyF4Cu4cmLXWCF4/F9Vc+iLhFQ8N/ybdprc1eEDdK
0KwWWGfYxoFzA17beqGfZg7dJUyXobXC0tPOKJURQlsj4wOdkbYJrdsA9Bja+gaGMZOMRBrJl6Js
tUHKqPM2lUU3eyXDxC91YozrmkYDoxfk3e8C3jI1b6BojT3p+OBholVOY8GsPUjHUV19n2B/cR6/
utQ2dF3TTXhQ6cEfb5HIKsjkXRBRGs9sv9+ynczHdU80IYOGe8bmgtS3nM6krdNomWCZ4Teh0MEC
AMi2a+09/HmpPLmleE3HDgFVsWTI1ddA42pTLDDqUshkeMNCloXrDvDj+SI8/UMJrdQXMtbCNzLU
t4K/b41MkTHBesTz4uDCmSljibtARXeVza+ewsS0pS7FR8e8t4nW/Y6Mdl2I+K2Tsh2lQKeXIC4k
xzCwMTM2uNmnv095Yh3TmD9quJzfFOu4j72mn5bz7Zal0bFPSj1TLFMOFz5XOdn5Ilur4pxrqw97
ORxvCUqyFvxg+gKZW5odnihwMtp+u3jAQr0QBFfBUZnaPEY8dEnwG74x6iGsNm8ypBtYhmNddfX9
CqQ7wYBxWhgL2Ex1kAP4Gu/18mMw7TOWFgdPCA7AhzgyqOl2O51rSS0UxFNYAE25KFtyXpDnVfp2
ES1WXYWVMQ641e1xDokDGzGdxgRoxO1yGZ4CGyw9/Aj14K7fYPc8PS7GCVVyelXP30fJu4m9Vyor
y5VrKUv6Fq3AsgovTy5edXXoLuRaQwoJ1Fds/C8wnzZ87fvaQlarcJIK87QR0QuK/rb21JNGVU01
OJybItpFEytzkMHzfTysLc2Z/nrDG4r6TRjR0UXNinkzf88yXdo1dJ/h2sBqcGStTc5FmQHhAf1O
AUpDuCURzEM6ApxbkshTxzN2aeR/R1n9RhSpXDqd082jwhcI56+dOuoFCXGWVV7O2aL9ok/4Js2G
jHzxgJBgXwKFSR5CPiobqrzrKYWqfSU0gOr6qW4gpx4vjnaUt/VeAefDfjj1X36Tdtfo1l9fmRsI
f5LWHh8TNZNtsMm40aWRDEG+D9Tzt4gi420YEvP3q6/UG4l6MByFpPkASP+kSzPiEi6RNItXDN/G
GYZ6MXp6TOK47zS7JEfHuwF224yJT4kBXbYQW+xadKLo0eOtfdbD2+I0DT/VVqyFA53Xo+vwM5Sx
8/HvKM+LazsjZFnhwMEhXKvnN802pAjIulWooWdScQU26VZ+zNy958RWBmahz9a9IK1YIqTwjCZH
tbHnshlXYEIz1ctYgZVkASoBg50WrFEpy65XZPXJuNcM49t2hQwFAoRY2370aO2QFstf+Zo8gmB0
g4egQrAVvBLszitpP+t3d9J2PPJNr3GVGd4y47vZi6u+iebx/Fy7CrYwj0jyPi3CcHXEmYAWSAvW
3WBEXDzaA89jyccfExgnaPqlqGnb456kx6bbW8ixaIU1UfvmxW0Xt1NgTUmja1O++CCqnJSp0Q0Q
WnFzrJFHzJJcdvVlYsdNX0E0tftBZ6+7qNWYd4XpWGLnPSk/HiT6XX3De7AYrnmmH/WwVZ3ub4UO
IlSU1hxmKiVlSP41zDR576pvqk1G97o8hlonX9LiGNNfEvfv0HA/NcVJgKfd4bq4m6jTmwV4RcvS
iwWsniZDvU5jdrqX+yNl4oQla9dK+Vp/vTTq0HGpr+yYGOLNvmIxRBJWkcc6S6VysjKK6jg1T3uV
/etU5LAsTuInn/CzKPzYp2koCuyQftNhsvG7YpHzSYdcDRNpMxXyTd144Na6lsH5xpFA6LZowTBL
stnVDQV9K/Z8QzvbCNRgRLacNe+qwpBgOL2WPusqyTiNLrbYR+3G5Ia2lSB7gQXEYOPCgABUV1FO
270z4c3s1AwIO6Y69ScIMxB7JrgAmdIAv3sj4l+mZjYZAOcmes8B/gfHFrkmW19Hq+ARO6p+z3rt
wRGlekcriII1z3vj4NX7ye2Nr2UNop+ijlWpPmECV5SafuQSXmOTBCzuw6+JXLcH4WgCx/wB6cVl
aFdKwe3yK/Lmbr9+TwDIJs1LExtiJmeet3dsvXiElX+A43MGPnhyVwQbbW4yYPHJwJMtlChfxng3
elZW7bkN7vBy3gvRdGWijRjMS78ub2hyv47L3sAuJQmz9gXGNIdybunMSfOj6Ir7EHUMmdDXVJyJ
swOxPTwVOWse80CoIuIeyyK+jflFAM2Cuhiz3TVHe3AA0Qho3MnmnOeAHbpusgLYPwub92EeLvyk
3eVtbmX6grBfkt07MhpTye4qeiDvoqrmL0fPbMjtgX0ytnpQWK/Hg4KDT5UZvdRN3lNhixsAgNbe
rNNLGWf6VL8ZiCYY7t5yqZy1BWg5OomE89lDN1VFTljCrWS38ficq1RfSkipv/oJquhrUn8zh1ty
lGC0NX6cvzpi5Nu12/F5hik3g4klpofCA7m7n70fjvBKJuPsbYoFbEDhyi77da+voSfBpB1dJdZu
Khb+R4tzLoy6bt7i+erbK1AeJ0WmkzyvnJiFxwK8mmbtNbQ4Gdfyfd/5We2fLZXGFkU9jOX/3Mnp
iNdj7M0eyMeS+5bEKp7YxZSxmtDqgZL7asqLsajfzGAG8qkhGN3m89AxVGo5+4BOhA2FEsMhgtFL
+d1+e4FI1K60sHpkPU6lU1PsTYuVnzKbs0imGJxsCcc542WpNwxUdiTN+z6yuwTGKsq5MCHI/UYA
pAawqWJNaaxG8txph3YUSZp6CDQzH+etmpTMdqYGjekJiKWn0kpqQpTic53a+cCGrt2HjRPGWnCn
ZlAS2tFdlFrBs45eJA==
`protect end_protected
