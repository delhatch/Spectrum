��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H���*�;��&��x�ʴ�m�LH0�A��PK�9��n�M�;��9���#]��8�܀u.�eb,P|}l(���πi�?��K�j�yؔ(m��_,'-��Зs�D���+�Yt۹�m~�u��t���-�O�@�
»�RY��5�O�ςv�/�-�qS�2A$(����vsΧ�P?��!�H��Յu}�[�C;L�o�!�e9��P�u��5s��H$e��
*�^[i��"e>�޻m��"q�=����I2�9u��@��:;/L?4ĄǦæ8}d3
?�-W���b��tx�j��:�J<�`l���͂��фV�u��A��}1 no�
³/a6[��!�ƹj���]dr���%E'���̣W�Cg�n��f�L����Z�P�:�syB���L�R�@�d�
�}҂ ��Mx\4�`0��͹ �	/(U�󃇻� b�׊�JX�|��9���	uz�k��fo�j@�#���<{_��G�$鮀��p�\��	<�&�?EPZ��'��!�uz}��jB��l! �#����%6�~+F��f_>�ZDT��GSYm�Tx{���8`f�����%�Q�c��V	��"�^P x�Yh�HV�l�]9���h!�n���Y���BNa���6���j�H�-䞹֓ե^�~�e�1O">��$�xv�.^S�Z;�S� ��M-�'�m_�����j��o��R�(��U�J����4엣���\ ��~^��7�XF��ߞa��G�	��
��nf`*�����N���|��` �E/�Y�^��Ze�90�Qz^�c�w�|�k�"��&�.�c��ߨ�[ة�_����fl2�C��6�4��J6@QQE� Ѫ�M��AT��p��n��"�Tf�!��e�"���*U����>�[��#�5n|�&?�N�V����B�+��Ȓ�8O ��:{��hE!����0�F����L�ߡ�%��-�y�J��#X���_s/�b�  �X�=3�N�T�P�O�5l�}H4P��W�)_� 'y(�����!8$й�o��1�0�����c���{�gW��7<��(vP�L���U���1��7T�,�����d�xD�j�1�S2�<�9��R y���BoE%��ԝK�O��n7�!���b
%�[��ή�_J��y���m�(�*R�e8b�=�r|
��g�#�fu��0Pv���t�P��K���ya}�NV?�F���D�d5A�+h������i�ˀnTJE��v�8;�
��`k&�a�s����}�}�w>���L�V�w9w{�9����;4��Gᇎޞ"��6������啼`�	�欫9�	{�ۚ32�*���FI>!Ƨ�&��d��YZV3]2A/:�n�3���S����JNb��8#�|�hGjoG)N�$"����'_Y�T����9�����rwl^!��M=ݱ��C�d�L�U��*�\BH���_ޭ�ԩܮ:k�Ƨg�z��%�L;�e�s�l
����x!��S[���	�t퀎�^x�VJ�p�X���~�Z��o��3��	c�������b���%Ú)R�J|���jG\@�z���3tFw��ĺ�<?&3q��@mIrernɧ�!�͕b�:���C�)�k&;oo8��{����ʽ{���S�����������RT1әH���h����t�.���E��DY]G�VS��$4�a
v���Lq���c�<����:7��b�(a�ba(��)�)�*m�Lt~IA\y���Y"�6��y�liy�<A��&j�xP�*EG��܆�G�d,��r���Z<'�di�?pᩄ���4�ī��AC�(ę?��ɦ�>�Fd�? �eR}�VB>-�$��v���W���$%��.�,,2O��w���FӨ�U����R�Dg�2���;�п�m�Z;������|7u� s.T��T�?r��=�J�c���ú���o�?bl}8��<��Kw���:�X��]��lf��6�P�4��8�(�C�q�
��˲W: !�6:�(*"B�55:k8�/����`��HG��UJ��������I��²s��W��F�v��E#N�0ܰOs6@��g�u�ĸ��w�)��"8? n�յ{9�㑸��ሬ����8����H��L��{Jsj���7�6��ɫ�)b	���`X��J���W����nE��k�����+��[xV�\��d���M� U���cdaE�!�f�������dfӾ#k�Xͩ"q"�h��ߤ��K\�砞�����o��]��o
%X�yu%�f�s &B�B4DD��*t��������s�8wحK��۬���kGj�k8s� ���u6��f�1��Gj6����2�M?���ۛ�����C�����E������?��m�n'�D�ɗF�@�>�J̴��(�H��W��H��^��~�Y�Cu��l)��D�L���;�0�L;��AlW�7Uʦ�C,ĊPv�"�X��Xh�'�����	A��x�M1�H"�"��*��2��	��^<mY[��y=��Ko�\rXtXP� �B��C���1Dl���2U����A	�{�G"�]�Q���v�d�]s��w����yϰ�8��2R���WF��%?,F�asc��ɶ���l�_B���M���|�aw� �0;Y=?m�cl�7~I�m��NA�������trif���QQ�6�_�-6Y;2�n��/��2�F�s��Q�Kb7�bN����pY�X�����c7U��>~�c�gC0����c/�d�e����a����)9���D�4�,��v�<h�ȜGc�}Ǝ�R�p�b  �	��@�RjAu�?���̚�aU�քF&�V믜r����{x��pz�(�d1����|�悀�Q�?`����Ҧ�W�ܻ<�(�����mɑ(��˷�kw�*��E��H,�;�ff�X�^����N��/��=D ��o3F��V RT���QLԍ.�y�#�)|�]t���be��X��OT���4��E��|�bc�|ԉ�O���'�W�:�A�� �9�,=�d�%� ����N8#� D��DhF�	��M�q���G�8b(6[��X�����!�,�ﯘ����B��5/p�q�xq��S�0!������o��p]���R(c�d\-�͡F�_O#`�u�mԝ<��f��8R�TE�r��%��0i�����0ƆS��؜+��YR:�ꡓ�B��������[孧)(B�R�nc��woWgxi���ѝw��/\�� �|�Y���C�&]Bh�.X����2u	v�!��-^U���Ⱥ�m��(ݺ��{-P��1ˌQ�+�ԇ���!�_A^��*hdA��5�n.��Ë ����w	V����MI�L�>;�U��f*������+P�җ����*ٮ���@�UW@�� &1�	~t�y�9Ўqubk�հ�[�;X��a������٦��)�8<�Ht|c	���6Y��9��i�	�mcT��h�"�@����7j��7���l;���~,?=[�d�-��)|Z�ݖ�UI�4.�(F��2���@�N�b�kЧ�H�K��B�&��I0<��)�C>�����CJ�J�⭅�������2����K�Ɯ��c3c�b�m������uH�����p�������A��,nI���!ͧ�BZ��*�t�<A6�D!��ʚ���Ct?n"l��3L�j/���}�Om&��ĉ�k�/��DAh��Έ$}�In�~	O������C��h��7��88�|�ك���ez#�Vף�xA�]d~\WW7�V�5���/�&Tx�\E��	����Z�u9q��a���.�_L��ǻt�#ar�]�̞q���)M$�
y����H�l��DW0�(]�<}�z������R���;�ɱO�/0ڈ�\�?���nр�L,D�e�S��B��n���"e~־��2�ltRVn6,Ӳ��χ(��� @����a~��h��ώkhe�*�������\B�]*�Vc���'���&�kBXd�|J��<_A��G�^%��Q���,m��x��v��~ 2H]�O5[�9��+�I��9:1�~��V{��\7������0�/��Pũ�����s�Н��L���$o��@pC�.,H|��n$���k�����I�/��9I2ՠ��Q�އ��Y���S����a�t�*�Q�_Yt�Mo-^�������/�1h���cx*���y{�p�@��<)�TR�F�ݗp��R
�M���=�z|��h]�Ǐr����f�f��3��3�/�+�a&�+΋�8H���*S�� �_��}0�(�E[����20S]�kq��P3�����n�ŹJ�VŅu��H��3��A��+�5�ShsWz#`6gt��$�y�"B�]�ئ�Iq�{Ԟm��6#´���MB�o�K_�jg:'B�4����v*I��n@����)�?��R�<q<��7��c��l&�l����"��A�hH[�JŗƯ�ӧ��i����� ��.I�VT�!�����Z����D�?h��UtZ��VC>>j�)ʋ����[���ݚ���h�3Q��hqʌ��{��i�P%a���AC8
3��T�B�c	Ͽ�� ��DY	��g5{b��'�� �7G��,�E[V�=���{p<�<��K�m�������A��83D�8|�_���g�0<r����9tU�kT;���>C�
l�~����'�ȸe�x���� ���[#�f�H�w�S�DPf&�xN{s9�]zH�Aɬ2u׍5 �儝�a�S' �^wh���ȋ窪螇�0��X�e�ӃI;U��r�ԙEg>Rn8"e{���թ!ʩ���vل���Y��c�v������L�
`O�:�BYiCwB>+y���~1��Qc4$����� �z���g5*I�Ǎ�	@���`�����N��&ׄ�9�����#�}�y,?�*e�?
%�8e.H�]F9�Ҿf�6�*�]Ȳ!= G6�<�B�-�n,�ߘY�00\����=^���x;s���C��<��D?����B�r�h:-ʐ�Fm	����>�"e���V;KG��6�V<3B[j(Dqa�QLi �A`tr�C�+Q�iL��(��L�1��_�MMg��8$�%f�'~;vS紑z��Sr����� ���M�N�$�mr<�
��6=�=����]��;�c�-�$�1��fUg�������R�!�5��$�C�^-j����L3�9��e��'K f[p}R�Y��Se1�����f��n0d�n�aʟ�<x^� �,o��R�(����Or�XX�Z��2�U�(jX{)Z��.����5��7��d�Z��"C£��'5H` x5�'Ǵ���uU<��E����{{\,5���I�.�=8W������n�@�R�h���*��1���5RKv���s�����=<�|1���,����(~�ஐ䳴����tw@}����w	�B�ȼ�~��%�_�$N��]�9���n�$@PP	�L��N�e����_ ��\*0�z��9×^:�X�#�t� ۈ�����x��oY��X�~�)��ӕ�o�{q�wp����1�|�g?C��N�G&Gc���d ��KN�W�T�~�0�%r�j��zj_�M[UDM�W`-�#��u���C�!~rn�@���Z���*��%1��D%�I�у�Q��r�%G��B����Es<f]�M�S�=Fѓ��dU���1�Mf��\�pR6�r�x�$�RZ����{f��}�0�0j��;u��뒫�Ƥ3p��"U5�@~hý^��	ۑ�������eړ�����Crsq|�����b��VK�t_�y�E4L�����2t1��o\�֨��(�E�H�'c�;����)��
	Q�
D�v���N[�cC���qe�㥩ήԭE9o�]�����e����|��Y�U��m�.���'ێl6
+.�m�W�'²�_h�tm����F����>��I��ⵋ֋9�"�dS`�{Q��Z�\i��"	޿��qN��E�^\K���"����~#�ɜ�V���Z�i�FH�Liq[ٯ��Ù��r�T:r�^�#Vԍ.7�<��BEޥ�X�!�n�P�M�JD~de����~�p.�>W����t�������� �O̦�9fo�Ja�[D��� ����Wδ�e�](K�w,拋�`6��(��h�{C��wr�����/t�|�m�.��)��S�[	s�KB�c��(���{�h�S�s��M>1���vO/l�e�g/pMq|�·iSƶ+.��C-i+�o��~Zm��~B��^;aHR����5cT�n�3����%�}�:vx�����)��+��y��-�Vt%1�ʛT{��*��C#�n�fɎ:!��^�Ӫ�<�>~�������y��>����
g׺�[ :w��r�����~y�V��Z4�w��oGEÐ�gdx@s�6��ۼ�(α��D��	�x#����'�{��9Ń�_Nk���>�+y'{7��(�O�BE��� }^C"�6�+7�d��%�d�*r@�폗�{^�.9�����L�B�Ky����t�Ĕ����o��j��L���`W���a(02�'��c��cuQ=@o~�����fv�xk���P�w:|]�R�*��\Y WGr�v���'��	����R�;Z}���!jU>(L��<�;�S�Xݴ�|
	��8��H������v�hr���=`�L�,Υ��:��3�wK2<S�y�K!�D3U���#Q��th0f���+�����b���G��]����L�r��թ}��N���@�G�FA���w'����v�]��$uY���-���k��o�<s��5):^T��U�P��wW ��P��3$pK�g䋎��|��ou�� ��֝�a]�0j<z����p�n���0�m���7*���1�����r^�����8�5@&2�%d.&�i

�w�W��W���`����~�ZE׷H��g;�ۀ�Ou�2���@�5e���7��Tj`��o��[m����4m�~`>GV�e��l0��p�6���:����ݜK�9�5�{���%P�A�FLp-&bKG�x�^վf���� ����plR��d��:c�[���S�K�m%!?m~�d�^gAyg��(X�b���i��^��\��PПXj�p��Em���3�������TF�l�ٟ8�MȻ��$ʛ4�<��'?U	��4T1 �2���|~�W�(|���J�@_����6�L �����u��*.�Yki,����ET�چ��z��;���Kk�ؕD�v�Vn���lqm��0�}��F��ߠo�#/���*�����^Յ|�xt���Ep�~b�(ߋ<��0��.~L�SS�mO���U|$;J�_u�,^�S�)Դ%�{���� X�,ݡ�����ɘ���c[b�,�Fl
����1]���y�E;,2D��9 � Ww��<X_;Kó�m��!-������@S3k9Y�߆�e"c��W�����K�@����/��%_d���	=�_r$hT��c�l�o��u���N�R�I���j���#�˦wE��#TbCD+i��[��RY�V�~kzH���S��ɐ�0��_-̓bGsԤ���{	f���G[���)��ԭ֊�W�s�%B�o�D�5��zl^h��j#(�5���{䚇��ެ���5��Ϸ��&�xm�tC񅊹�ыT�>d��Q��!�*�L�Ń�21����������<��+m.ݺ�&X�k'ף����?�d�)�?�P��Ս^]f�v�?I��Â���A�E|�5Ы��uS��o_A�"D�%��R�q��9��e�&��%B�qjh��e������x����G��w�_fx�>�Kx0����@f@���b�>w]�Ǔ�3A�Y\sc�>>A�>�4��[���ƥ?]/x�������Y ��Uf�H)�3�ٴo^,8�\~#�2�/��A!<��(�^���"1u���J:�IFYR�?졐S��oXY$�s��M�ퟦ9��*��MC	���Hw� ��-�-=�����Ms�)����8q���o	�@u$���Ɩ��53gZ��6���<olW��r��&FcJ�/ux���XoH�BG�[~�->.�#Ln0=Z�c�\l.򧸬(�v�n���󝥷���B5��SW�i,�Ōs�,�t�$zx��5ǪS�|�,����8���W1;o@��N��Z&U-y�+	G8�F�w$(&�������~)��jq�d��uT1�ڑj�Ħ5��aa�^H달�T��
\�����敵Wk���ƎݳN_}r?o��>���J���{����4ɽ�����4���3�`=~1G�-]��󃹺7"��M���쏾%Y���ߡ���N��y��h=�W����qFv�#��}�j��,�I�!�����$�[�xⓂ6.�B�]�#g!�#;_�i�]�
{��bF	��=�L#f���U�j:47q�N}9�n�.1�y�箑��:�4O|q��;XI֔�G��R��x=Oc6գj��!�u�(L��ӂ�(���������u[��`���y�_g&���9���_�}�_xf�/�(U��.���o������v+m��9~E�$�D�<���S-�����]�%,.9P��R� `��"e�>��q�r 2��t��oh��,$O�n���0a��vA��r�Y�<�����
��yԼ@<(��{��
vݢʺa)^9*�����!k�x~��ZT [x�'��x=[n6��1P��c�N�ޞp��"��$=�s����xnwF�9D���;?�Vw��tg����#з�x���<�N]e��"��q_�6�°\xs�Fe��C��D��/�T�y�Dp�+ �w�td� ��Հ�7��֍�(�D �Y��x_U��ݪ'���%eSH�&�i��!��ӿ�(� ��j����%����=J>d� ߎe�?�S���T	�'��ŬW���?M���4�'L&C��~)�'(�$�U�=��SH1�U��-7�%})�GLgk"���r����y��P@��_�P�3ʫ���Į���t���yC��CM2Di������zz�[�rwsl� Q��>�Y`�?ԆF�{G��fS�z&P<���S����^���f�^��_��$g���<7�����۰������W���qK��8瓕�b=�W���j��7�<)���
���(W�k*�)���	I���;���pl{�	�?,����l�*O
%�K�⸌i��.'�0^�]�D�>E-5bT��~Ҙ��S�-[�t=l�E��U�'����Qk�d��]�)��H�?�y,�2�I9�����vQÅ$��<W�6�"^%9��8���G砞a�"�x�Wj��Js��)z�F��ZP�,ໂ\������%6�s��h$�]Y���"<+ {�\� � "��Y)b�������T�6p��c絏����JU�� �ҚmG���
5^���FʮV��wֱ����)�h�
����E������09LS��)�>��ܬ&"����i�1����1�E��,�}X�1���e2��!���q�C�?��qi�l�����_�B>to��gy�ʘH��o\�0�y�χф��n���
�փ�]濩cЛR<0��U��ko��<l��q4h<�D`^m��Ԕi�����X�f�)'o%�Z�eμkW���ם$"B�|XWX��k��(��Zt���x h��A�*(�}��b۴!O�ۆ�xp��8��^�!<q�,��)�ϊ����
��Y�2fV/T�-�+C��V=�l�0$���� ��E�-m%�F���i����8+��C�a������f��_g3��6��H�.��k�7eBM�rm���<<d��^�CLLh�NN�0�m32����h���J��T�\7G�~۞�^'���SD����L+��`ơ*�f�@�)$"7�W��-��9���F5)��a�D'[!�}U$66ēT{��_��,J
U)"�t�\��|�1����Q��"p��B_�;��׎%q��APF�[�(�?~��,<!CS<�/3��<}\��6P��mwP_ʩw\�����#1,�M�1�(Ad܉�`A"\��|w$����g�]ϭ��-��YP>V��R���	��Gs��`�jdR�G�?^�w�(���?w{1���m������%]�Ei'��[+"�D��se�(��a��*���D�;�HU�9��rލ�a�(���	�G98D����=���H��,'��	� <��.b�BJt�⇏�'��D8����e�x�ΎzF�v�O#F�F�qXc�%0��9��Q���ey)�	�By5(ߪ�ȮO��@8O�MC�y߮P�c�y���U:	[������l������n�	4���՝"gߠl��t��.o*�^�l����7n
��Q�.�=w2���q*�*@�Db�mԠ�XWf���T�� �f2Q�\N^�O1�$��A"�1�^�P�sZ�h\�ZLV�L��[��fr�M�%j�lW	��H-�� �%�p���˨����i����ܔ~�����O�j숬
S�2��M(��tQ�>��<�*���H����`]�DeM|����0�R�i��z�re	G5����dg0�R5� �.��?��oK�2> �/z��&y60vN�c�t,70��H��\�XV���(:@*���ݔ�N��8���J������e%Za�R��>&�3�k���\�\�X<�t|] F��#����DH����p"wY$�9`�\�P�-[�W����*H�MRԊ��w�g�w�'�w�a�z��^��+����/cc���ˤ�m� n9*��g���x�I����vZ�j��5��tuG�����ԛ2o�G��p�)6���N� ��������?��������j�8y��1i�g�H[�� r��N��,�&Z�g�[ȎS�1�.���n�Yh%�vEb!v%һ����cn"I3r�W��a:���"�s��Z���^�8"���C���o���4��*�JL�5��R8�;ki[�K��{������P�R8�.83�=���2V�iyg1����w���������F�8�^}�J�nJ��`�����bh^�r�0���(�c���2JBEBפ9@���k�SO�d$,-:d�I,Xlo���.S��l�;�S�+)�d�:������]vjd��/�K8�p�*ۧn�X�C;\�4�Gm�NW%S��&��h�����?P����&ʭ�������+2鑓�i�x ��	�	6�̚C�xk4=�r�X~�^���M��yS��mC-�a $ !?�inLa�P5�ܿ\�U{n�Y�+V��R���kq��;*�#6�&O#�6�_�0��Q�剛�x�����?��b��GfP�vmCo�V�����v2B4�~/f�T��&z�Y^��v�-��W�S.�(�]��M�X��M!�o!P��+
R���|Ek�����?�Y$�äL┴��Y�gвE�0��X�`�Usy|�NA��4�t��3�g����3��a<��,���4]�����v��~^t�RuiՌ���/1�dAB|���CR�;M�*}�%�d�9U
?8���{��4�G?���tDM�������ٳE���{Dv6��	�p�L�ք�ߣ���=g}��U��P��X�9f�h����@x�����l�c�9[kb�/�=�����m#3��v��K�$?k/�v��jJ=�r���R`f���;
�!	�Cv���V������,����x�=:���v�j.C�?���1U~�ƀ�;۰�	�5��C����2Ⱥ�o�f��j�����|D�'Vѽ.�����-@����#��z�ւ���9���6�a�#�yZ!})O|9��,����������n{z� �(��!acZ-N�`��$�Z@�=�X� `T:Rmxp�8=�&�sa�XQ
������w�6���)��{�2f���|�$G�`�]ʊtR�dj�V��>��`C�2V�����n �9��1٩�1�k:�"�B��Px^	��ע&PO"d��A�	�jL�Aۄn�{B�dZ�oc3����n[�x!�jw�f
6a�������E�Y@$ ���7AXnbo&I2��R�6j��2Qg$䌐i�h�yr��
��b�N�dH�"Tr���V6�23ԗz[X� I���J1���Bx����u���k� A2A��7�Hv�2�0�G���'���k��=���X{�:~:�f[���>�2�����Y}K��L��}��˯�t+������ŝT
Ik�1�����HM�d"'?.f��e>�qa%�cx9���ㅢ�$W@y3�'��I����w3�&Dh{����o*k$��kM�����/�L!�7[��5"����+mM�)�}X��k��E�=Q�n>���w���Zӱ5e��8�oq(����s%j�S
^>�\�OFZr�.��R_'i(�m�C�(F��F*�p����Ң��o��p*�+�ԅ�Q9��q��Y$��j go�1�.ؗ%@�����>���ª����'�)�y�26�W�D�Uͩ��ҡ��,�Y�<��L�� nCt�K;n6LvU����>^ϐ�1����`Q1�nvK�"�iW��d�%F��J�X~6y�N)�5r������.y�w�G�R�L=�����?a�T��;��%����֒N1s�_�r�M*��h�- k��Y�Ѹ�6��.�㌲h���[\�v.{E�,��Ѩ�g�֩&آL^�q"��]�>"0|N�C�����iRq ��t��@�T!L�K��	[2�y��=O����:&B�����i�����ˍ#�r��o��%M	H�����}�8��O�io5�:-ւc�R��u�A�[�.�.c!V�1o�(�p��b��W5h~��(-]�y2��hc4�`#��@u���dS�Hv�����8�Z7�9�F �����d��h{�02J6��j�+��TÙ����W�lc���cǪ{�PH���Zf�p��Ea�Cu %(�k��z�:�����Z������2A^ ,1��q�:���*R!�u��k��'���Z<FP��t�]W7���T��l,����!�A_��,�Ӵ�a���R����~)�BcO{k�+�xj��a̢_����l%갣����߅u���M�:N�����"�N|���š�*I{"Q�y&b��[կ�͎"��7Kv�.��K��R:z�0X ,[���k-~�7ٶ�S�\��k��� |��@�\L�aj7�ԉz�H�C��n�~�'��-nw{I�Uu:�`Zho%b�0�@
��WH�"-�����0j��otQ��m̕b>̂��ڙ�����^ߦ�h��%�� @`�@�?:���4�	���������y"=�j-����j��fq�U��[���T%ad{�,�����p���u1\"�Q�Zr�u�C�9�1r�!;Ck�����}s�n+��n���,ݜ[u�}*=D�9 i����J3�{��y�&ũ�Nn7A�a�t����/�nc?���BZR,���0F�rd�]�͇�[uw�����'���!�R��,�\Z%�z .����Ż�S�m�<���bF����O�m�L���䖻�$�y�.hH	c��-�R),��^�*)J

2�#t��͎vk�D�(1@�u=��v�<�Xc��)�q^<n)@���ǳ��=�
�G�f����y��k��-=y;��,r�N�c�u�ߧt�iȅ&�b:=�#�	k&r�<�39X灾y`X�z:2���S���-��I=�e*T�`;�E-y3�5� X��^(��R�>���Bi�/�^ �hbu��"��6�{ƹo/b��]�}��d����h!6 �u�{�m*��Ќ����\�&P��Y�	DHg~��9��b�J�\v���p#�_�6h	]\R��z�ߜ���R�I�T�l��o���x���ݰ��tp2kF�����c�T��g'��S��F�|��`V蔝_1c�c����BG���`\�2ZQ�w�$���^��۽H��g�#F���pl�˛=
��J?��u��έ@�n���O��J7�GK���-��r���Y�	�D����b��s��f}RK ��r�zƶg�@�����b5�:���K(���H,UQg���{�C�4�%�ss�Y�)M	��WR��nm�G�m�\�"/��ј�
p����w���,Q.���{��v�R��G˕��o�oµ�!R�u�r���C���/;��f֚���|;Bh>w1�ߥV��Nak��NNs[����#������Ћ��i�I�a�9?ܩ�����2���z�"��y�ђ�#[��h[�%�6�:���% +[���<@)H��D�c�w)���>+h�?H���(�U�Q��V(���9W�W�sQ���$ZA��C�W2A5D\"?�y�4�B���i�.�e<J���V)��
P;�1��� iZ���ؼbǹ�^�dsL���VV�[̲k���K�;�?L�6�A������(�z�_s��nX�@(@���ŢYհk���U4���&�ɻ:��}�z���2�<'&�k�L���W�_pT���NaS�DL�~TIL�aH����r�Grst�>�,���D9�'zWRj��+��Ms4������+� �L%���Dv�� tթٿ!|A����	�i�
s��9�q�I���m���1���0
�^�_N��/����	�7y&�)y��� ������_�zN�D��V�Rg�d�H�f��\��>d�W��v]� Z����[�p��p�:^�Tz5}Cu�YY���Ħv���3b�PC�/�G1�/`ړS�1m~��	:m�g�ĆNiq�B�s��ҩ��5Pbf�cO�ꖌfS~�Q9撚�?H��U��� ;ȴځۚ�*�E�<
e��3�F:
��F��s�,�n"߹��tEW�j��b���H	�xT�{4�����q0d���
3T�"�-��p�X6��3B�^ڶ^6.3^ bdΝ��YW��U��p1�N��D�K�R:Zw<�!��S�)c]׼{�(�b���l2���:OŵC������JfJ����`/Mo/����F�T�Fc���'��s�?�g�&�)�pW��%���/$1�tO���0uC�w�t� �rÁȞ��j�N���\μ�)��S��Rbz:{v�ȸ�B�;�S��x-	������g�&��yyCU�1�C�cƆ�G\��b ˛81��6�y��ѳV�q:Y��z�P<�U�޲B	\Oc�X���x=�a��.�=�L������խ|��6X&*mS�x��t��Nt�3�Ґ1rv e����]�Ez�T�V�ڪ�A��-!5f�=h��W�y&)���"�%�CBY;׊c$������CI�1{xO��m�Z��!��ܤF%����z�Φ@�Q|ށ��)5�[j��:H
����R~�o��W:�}QZ�k_�{��ᝬUꢄd��7��gH�D?��2���m��c����X{�[�#A'�?�\$?�΢q�:��3����	21Ȅ���esb�&	��8g���ۆ'��=̼i�%�MEa�A��Q�S�J���\�qy� ߸���Ue�L���ണ�$��W,�,�0l�J��� �e<	�{`��Jy�mc�f�7S���x��D �ٶ'��DwF�9IlBm����UG[F*v����26bt��Z�7��y������}�L�"����&"����dm��!U*jm!i�|�-��2��}����#�oɼ���S��p4��� {ۅ�gE�}���2D�B���O8��l�ۋ�3D�}g���9@\}�>�"����VI�:
&R _P�^-�讻�T��NB��e*.��Hh�ۣ��Oo�h�Ƿ9u�@/?Ժ	�����?�47V{�zLQ3NgQ�2s(.��?�e��M9��)ML�|����wM�>Z��>���Z1����\�W���F�7<'lH�%�a�B��q���X��b���4=0Wx��"F��Y�� ��Y�	n���p; ����G}�#zJ ��ʼ��+�*�4�ҙM���iLբ5B��g�eA�D$VE2��U��@�B�t�z���q��-b>|{�+�	�*:Zս�~½͆;�� yEK��j[Ͼ�N�-[hKiw�Z��ל����)�>�d�b�@Ho�����A�}�S�NV�t�:
�k%G��`o���uŻ2VyUܛ���B�d�q��0չ|n��T�H��Į��V�u�x��*űRw�<�I���8w޶Ȩc��omm	)� �2�ɧ���Ɂ���5��J�-E_s���Q�T�i����u���0
�x\*[]��ڨ1�U�c��E 7���vt�`�:��r��#t�t7��	�bh�"�T��oA䒑�_��*� ׺gŒ�h@qY��u`�hY+A��y����PF�T�R�ֱn��^�š��1B�=d�F����k�-�uP�2L��¾p�Ya�KZޮ���e<(�d���ƅ�|ad�tH���k޳��,{���:Ƙ~���kf�%÷a.�����U�b��X��ܙK�w��Z
Qږ���5�E4�����\��F��>�Xu�(+7���a�O��C�i�sa����.��:V���2�1�����Z�޻AJ��w5}��m�C�;�Hn��qD��[��x⅖�t^����&�PǓ�wU���Վ���:�&�'��Y$�wz,?9<;�$S�l��ʇ�$��	�1
�T�.N��MX�R�]Yj�9��d��1@@�R<�f����pv2�J/][����]X��y`�\�e��q�D��\:#[�q����4��|��55U
(IP���k�F��>�T�|+�W����i�&AM�h-F39�TG��� aq�*= 6�9���ȳ6{~?�<o���NO ��h��̳�\��v�̦�e�����m��.�"u��5�#�L�D{9��8�ւb������AK��]%<'6��7O0�'�FAM���t�����l)��8<V��r�ao�Op�1�.�L+�A3�[��F�jͭ)�`b�b�\/�C�Ŭξ���e٬��ن��tc�5��EO.�([��>僲tޝ�}1%ԇ}�^+
e>/zB��,�Ȫ�yJa�2E�q�	�,�)������S���ҰkU4�jX�	�q�,b�s�V��edKQ�s�\�=��m���\Q�Շ����n�ON*����>K�6}#ߑ��u�TO�[��D&�PR�]T[_�'�C�,�K8/S�g�]��f����}���$�$!����%���1G&��]��g��d���K&����A��LT6˵���aӖI�"0S�ġ�6���8c�Nx�<[����ZDNd�T�3u�?@q�Y@��xS֪��p��O���ɩ�RU�����bT>6&x��F�<�2������|��7*�+d�t�eLڟ�a���-��G�������O �gF"����ɄL�k�xU�{a1j
�t6�9s�z$�����T׈6���!�lI���`��1p�~S3���)����	v$$�e!�	)!$�/�^.�VdV���;���dӈM�G�ʉ�'2��|��� �O�z�u2��J��A=:ǎ�|ܞ:�R�����e�1�I�EjrL���&���%8Ҝ�C�-~�yd���@�i=��t>hy�Im��L$'v����<�%�oFyNK�'}tHq�'�o�^��l��/׌%�ORЩtc���ɶ43��$!G}W���Fz[���N���B�S}w	:��d������Ă����d ё��Φ/�X�D+,��%
0����G:/=���('!%����&��P9��;�Cf�l��`�C3��;��G��x�Š�m��ʹc��x�0�f9l��{�Dzl�7�E��&��ʏ�Agc���">���d�����T��� ��p���c���0����]F.��)��_���Q�Ot��]����RYj���]��Wu���O����璁�����(?�鿛-�0�ϡ~��I3�]Rk��jq��׶;��{��R~a�޵a'��������'�p�w����^ʾ�t�J�(,�t���6��(�`Ң���	�ˎtbI ���у9��ǅRQ!C��3��9��[��&�ԽX�T`Dv@B�rq�I�̅�]{��C�/}}�M7k�B��P;�2S�N34	zA�(jSm�����/ͧ=��%/��mF��O�'#�E��8�����D����,6�Ky�P����7��0Hs�����5���x��"2je�˨�������P��hm`�JNV�i�@ ¹%���(thB^{����9�O�������9����r]����Qj��N�M�*ǕD�(��)�7tŝ4m�?
7�<��N��L;0n�����S�#��Wn�-�q���%�|�j#m#���F>�(��q�Y?�j��^j�UJoZ+H9h�5��`�w#�7Xw/og�E�9d+=^q!6mk���a�3(-1��A��wF[ �NI:%���h|�~���Clr}��b��:���Q����\8�Q	(rgI>�n�Z_�vz2l�$�����^�,i*��\�IG׉������M���7��Ɖ,z-KR
N�j�=���;-��~f��D��9����G���)�:�	����~ؤ�����,�5���C��Mc���؟~+ن�"��[��f� >�ń���PSZ�`�ڸ�C�fZ�`/��Ð��i�_��E�c���a��f
�yZ��I��v��|������o��/�^��p5����0eVE�&�W��;���U9 �_�Bnz;��]�#����u�����g'�T�����8~��>ܛ"������3"���u�\v�Y��� �����^�_���r�����pD�2�(b{��r�TR���珯��M��crT�#3d+)�O����H24ё8X�!s��}}�l���'�N>dI�G�4�%��3T��4�oJįv/�2����	1�������>�Y=��#N;������,��3Vg��U9�/}:�;�D{�GnX��ѓ�����,x��ߙ�O'b�W�V:��WI���#�1��4�y���z��V/��(D��Wr7#��r��A��lڇ�����-7N��v���E�l�e�����E7X�keI�w"�?'%���9m�oSn�
�KgG�W�Z��X�@V+[Q��;����"�~5�ύgv��}�
p��]���JNr�/���d���Z�C-C��a��"�W����/�(��g�~C1�a���Y)�q失��<� �'P��$�þ-�� ��e���,L�`+˺/�&s�����h C7��O�=И��h�.Y��#%�$z�\8ځ��#BY���ь��׮ǃ�{Y�e�^��`Wi�ƦϽ�tĺ��{eAB�~���z_<#mN�,���~�t]����J�ɸ�\����N�C\��%Z�'6A����(X��u�X�ux
�T�2j��-^��)��X�p��}�:?s�c1�,@��4�v�s�jl�u�������1��T�b� ~f��$�oNq�4pI��*Q_������ȚaI�Ig��x;
͵�
�*��*?�!%�����4�Z�1�U�F��1�p�4\W��#4ӊ`���0^��g���J�l\)#�����g����{�������vwd��`m�o���*��K`��{.R;��׮a����P*�-�����c3!����Q<جy���|�`pF䎷��C��La��ǽ�8a�I��6A*p���.���p�N��0���Y��]L��
�������_�F��|rlȲ{�+ȏ�}@e7�ֆ��$X��]F˙[P*L����k�QV�Y-�A[)��]W��;鍂�A�sEv6%����ӷ�b�W]�Z�
fA�{�)z�0%�����I����M��Q�� ��z�L�U(�+�=�Ō��V��T�=�
� �Zκ��D�_Q�4�r���k�`����r�X_�XLܛ�`Ū��h�\3�#����5����L0.6\��j�mH��v,fA[6q�F���V�w�e&��
��\�X����?��$
}@̽���aV�����ӽȯbARj�K'F�e��������$����gEL�_�>���3�sS��x��X���t_4]&��yF�iI�&������&,�9��3ӚA��KS�B^H�*��)�;�!��S0�rΒ#�/�"P�/m�d�X�tR'�7�hJ y�@ka�wɑ��%��)n�{Ĥ%�5n�T8�RY��T�⃥�-�\|����+������JP2�y�����m�$-tQ���wdqU���*|D^�����@t�z���X�U��O⾹UE�3��!q��f1�[��t�g���lT�ִ�\����N�70�i#7��!�P��h�x�r%m�c+�N�Ί�A�'}��(#�+M :I��_f�s���L����C���$\u�s�� o ��/a2M����-�����@�#�@#� j�;�Ţ�h0,/��%�`�Ə\9:�͢x�E>���~���T4h��72>��R�%1\AE��TRi���Z��M6�k��Pq:�6OH�����-|�	����`�ėV2���`�x@��֮�I���Y� �����q�ʔ,�q
N�Z�H��X{�2 ��Ͽ��P����?Oc��w��I�^c&���O��4'�p�~R:s�Y�b�8ۊ��^��!v�J+X�|�Y��t�f��w�{�*]�fg�w	_�j�B;@�,�U�Ʃ"�iS�c$���$��H
ME�ޭ�F�1�>�AgI�c�!kI?�g�ۍ-񧙎���W7m.�Ŀ>tlڮ�T94*����j�K����+��7?�.���yd��1x�PӾ�Ѿ��m5O���Ud_�L�fǅ��2,�.4�T�Zd/9f���}+,�p��/^#�ҌaQ��8�8���Yf2]�c- O�a6��w�;3в�yJO��� �p9X��|D�	9d��K��:��d�c0C�·�Y˥i�>���������6�(h8����}�)-M��3����-ˈ40��������G]h7$��XB�R~|���t@���:4��2�.j���RE)2Q��u枕&���'�"���'�ALi1^]n�= x��9V��0%�X���cIe�J�3}d%3�{�cF��F��12�ȼ�##����2�3�k{T�a���A�����#��k�pt����DITe,�����R̼��]w�����#i��&y.	(��϶r|LL���|�5�<���hu��bHD��k����F�OK9��_Tn(=�&���Q#*K�,�L�a��w�+�=%ig��U2/J�����+�A6�j*�0�d�!�;�$;+�-�BĬ{�	L؟���/+ǁ7��L��ut9���jZ�o
t4��?ͦ8k@�
�"���bЙ�\����������.��t�4(F=$��n��E�W>�Sҝ��%v�_�>n�3}鈍���3��.�[M����u�5��kCR�'V�M�<�^E2N�`\��#������r�#M�j�!7�4
L��F��b��y4� ���$��1IS*
�/�ݵ��nԺ�ʍR��_��2��DT�U+^��`��K,c�F�.���EY�?Ѕu_e>�`��ː�u�� 	N�ယ��un�iRJ���M���Ni��W˄� ��K�@˴�l�g�p4Ѕ�}jQ���u���R#d�R���%rajum��p�B���	�Q:jY�N�u ��#�R��Se�Ok��u`&Dy��P�M*m��-c5${l�~N��}��wj���3�͐=��gs�E�\�Y=`��[�S���A�g��^S�C�� �Ѱ�����Qp�LE/��	�^7d���Һ����)��@�{%�T{����{
�/�u�����6 ���G�����3��py���Y�0-��;ǗD�~$�B�!��o)<+sh��aʰ��A�w�4x$S���Z�e���Bu�@���j�&���R�/��x�Q��U���!��3�,�<���q�G��O��]��%N��'�k�{��<��8��z� z�K"����%kC�/�ץ?��_m94���G�<�J��;�ԅ|�����4��>z���N�˙�e9����˳�/�!4��6 �����U�� W�v���i�j�M��}3P��x���=����Ld�������B�4G���Ε��T�jR֠D,�ß� ��?J�*,`�֌���%WE�5����KXI0��7�:,�a/�$5Y%�@�RMa�Jcj�	�����.����4Y�qړ$.���K�y|G���P�YWb�2\cd��B���Jj8�/V��:��T��-�����3�m�U�[����˃�=���@�*4��]�sI��J&J��l���v������w�(��yRQ�[^
�_�&�>��c�C�>jԍ;�P9��E��s^�P�Tn%%�OA�x� P^칬b"=O��}{	�Oc� zI0��P~��`ma�Z�K.���$��҇�J�,���+F,!��T!X4j`[���#�E��)�z��f���ҏ�7�K�%"Q�E��u��1������'���l��/��c�{K�� ]��v����-�J�6��n9G��*�X]�'��f:��U��Z��-�-��V���h���k��+���2W���i���`E:��x���v��A7H6ҙw*������a��� A-�^܉��� yV�	v�g��# Ѻ��ɧv,�᠝a����W9��x,��,���X���	��0�52z;��0��l�J�,W<\m�R�s�������6���XtR&|r�Gh4FY��+V,�4���0�x
�=f	.�� wY��[[#^����w���P�n�s�m_�b���@ɽ��T{�Q�']1s�P�@�����S�J^��_�	��FX�ã?������'(��
�:e�Z�f�+�HGI�`�^RU�o05�Sw�-�u�X-df;���:��ntb�Ŏ����Hg�WpZ��ù`�;<zb�sr���Z�]&�Tm�����uQ9WA�7��+%��9�s�,�$nj�뜇��P_k��ơ\���>��}ag�`�Na|�8e/�|%�|���b�mPE�����iуi�}̍���ݭ�٢2<[$����9cHм=��W��O��G:WC
��?цw��W�	#�g�S��W���{�V4o���z] IL)���3QN^�!���X���qy�����O�N�1�"���N
��t�IzI]�� ���3�Ѭ8e���/y��KQΨ��: ��Ɓ��&V8�S���������ͱ���>4B6����l9����*b_�Ncm���{w�B������f�
[W�<`͏� )��gެU���}C##;�#��6�|�&�Z��: j7[>���wm��O!�S,A�\\�гҌ��p�{ާJ��U݊���,�Y�3]GL��ȯ|�<�KI� &�EK���$�F5��Y2(q�-��"�5�ե�����7�̷84�k��XGh�L�bTL7�� M���V��[�.�u��g�\y����-͋�}y�nǛ❵	C��x����F^���l����1���2X���j�an�a��䊪]�M�����#O��Л ���ir�ϚT�@��K�E\�e����:�=�z>F*j)OP�����$BȮ�N �A�J��XQ�,��V/i�P<r�7���Sg+	���s�<�ƌ[��aP���Ӝ�!�vJH:��	cN���\�:�&J�	�� ��䨩�
,��_h��  ש���ĄEa�#i���q]^{ꈀ�d��b���ن!��C$��d,�o6)��m��|bP�)�ql�y��|� e�)�>��ݷ�N���c��m�<�1/~ў�t3��4�Pg�t�����i/��r�gˢ>(&�H��2ܬEU_Q`�g����m�N�o��j2������~|��脷�J_]��A�BG��@	��q=ǙJ��A�X��#"��2�8H�(l'�n�Ğ�~+���!N���n�B����e��H@�$���R�UZI:���;���8|J�7⯱^�b�����.>ĝ�k�G�\�\�L������[d)@z�@_�~��,	x~��(R�A�z���r�����PMJ7��ud�Vᇡ�K������������ar1��7����K(���3o�i)~o����4�z�e��>��uD��wݭ�f�� ��b���(�yndBv~Y}�1YU����:j����b8ziK-����.@̖>8��q�+�ׇЋ�C��*�wNB8�!��E�ƃ�[p�<�1Ψi&,V�� �\5�A��y��Bz�iQ��P�wp��q�������E�K������/Z�M��� �������4�'�]%"gZ���J�r���h��G^s���۠gGJ�K��<�J5�;���^�"�a��4�x��):�k%���aPP�o�;�!K�"�i3�4-�2 g
�Q奤�����kw_���M܍-�?Rv��^w�~���.W�/Z�����x6�&���?�ۘ��UF!T$:�8]4�L�E�0�T�'�=U�9�����?����b�=X�n�[�`6s	� e�p*�?A�ﱾR���M��jd�ao���*D���ȋ�j��'�2h��D<]:��y�5��#�Nj誱��ֺS=Ř2R*9�l�lge`��a�6��Ö�'�yܜHc�,���H4�Qgm�g�#T�U�(`w67Ȃ}]����2���w:�!�3Q��%�(G�-�Ë��lK���{su���F�2�X׮�|�pMu���;s�&H�j�1��$�Ź�>�>�}�Сo��A�!��
�e�VQݷ�#x�D�Ξz�/4���>�5�{� ������ �������/ձ��b� y�_<�h�D�ɞ"_��s/f���{Q�7�ߝ�[b�E�[66]��L�匇.��0�R�(��gr��1�#�JC�E�?6�~̻{���������n&3y��p��F�V0�w Lj�1�\g�Ip4�aJ�l�����8Re�gظp��MB�.�t^0�&}�8o�̈Ҭ��5\.��W��S�P�y
�ګ��;<_��R�˨�ŧ N�av'u�Pq�
0�X�����^�H�������r��D5�Ǫ���!����-��)k�R���F,`�-�ԡ" O�(�"���MP[EЎ\&�92�M+��iRB�+��̓(E��u�ާ��Dp
�_��H0C���n���n"_��>zeN���nc��n����t�P���NNCY���,�3���,P���<��	��������	_d�)���bB
H���{e��_aW�z4�,�p�z��Yxb��@�|�f/�,�,`}q,�dS�O����������w�L��u��;v�d�V��&��4�{I�L8�g��?՞L�DF�'�^ɨyP�RGÇUn�y�Ƹ:�GG4!c���H4AM�1#���/�P������x�MDg��{�͝ka5^佟�U�C�`��h�//��S�OjJQ���F
�W����WL��
G\C"뚉���Y��$�tuQ�dV�Ɖ=Y�N���Gw� �tf�a�Ҏ�N�w� {e@i��w��UPL�5�Z�%G����n#4�$0����p��Y���<�d%y�j��țj��q%��ۮ1�����bց�abdD���G��A�����F���\z�Ǩ�u ����a����DU�f�K?��h���qi�j�$#�����E�� E-� �6�<�v�I�ݸ1|�x���uxm��g�;'�m�Q#T����n��K�@�P��=�Z$�q8ӯ�����a:�f�?��:g~E����U�=��6�)�ѼnS6�lv�I�����+�(����1�؝ 3=�Թ�gXc�y>���z��u�m�`�F~	$/��R~��UA �"�B�=f���a�Ygl��% s9y&��R���9BH�D���A&e�#�a��0/3�H0XP���ն�P��F��ga��w���&g���G����fȧR���;������})Ih:��^�Lb�sB�cT�v�3C:>	)�M���Yĵ�c�e�&�a��$���2�dϗ�+�o�b4���ـ������hm�p�@�L���H3n��mD�M��A�Eq���5*H�*����˷ikb�zC�V�1�y�d�p��Q��C;���:�G�1Vs/9�,�װ����}un���9�d!tS ��@�Y��1)m+�ɾ�z	��"Ѯ��n�ZI�HǅY%h	�~�������BK��#p������t���)�&��f΂�At����pIه�#��Y;�I��l�YTsuE��2j�6jB
�Fh�����(H���xeM�7�r�T|����VF?���Y�w~�J�I�x���$�+8��>9��Ϙ���;@�HRGPyh[��� C�Z�QS.؏{<����.���!�{3����ǽ��\s_F�f"i�n�����2�$&��Xp�>{�J����A��୼?	v�������f��#�u����4>�hݪF��A�Lx�4j����H��]�a�.��L�"$����UNsB:��sW\3wޢʖ�ְ��]n��`�o�r�1g�>=�>�J�gm��@}�<�e�=YC��*��o��A��������x�[���þ�q��$hi�ƕs�/�Ш&
?���ݐ�a�ʲ,i�������ts�n�o�C�S,��%L�,��	A���KR�e	�_�/�6��=ڱ�.,%}c��U��uخ3f���曭�"L2Y���9A�ۏ���i5�TD:�I�S�A��r��H�|���dVy9��9bi,ū�7�?�m�G�2�� -�y7�LTۼ m�sH(�W�v0tb�� @"�X�	����$�,�Js��/��c���� �-�=����0D	� ¼F*�Z�i�?��Ń��0z}��Dj	so�ȣ�����Pݪv�`�6�ӎ�R��R/�q�(�Y�R��se"&!��	�Z��-n8�^����Ҹ/K��I�2i�� mNv��˼,�[����O��3�51T`�X�D���&SAi!m�d���۸,$�Պ�4ҭ��~:�:C)��-ڏ����skK���|!����2N�f<\(^SA�$x��oW!��E�u��}�+%�܎c)ƗV�f��M.�㽧�2ԒRw��x�̶X`�z����˶;aK�ܕ١���vέ=���[���B�`h�Ǉ�BSLT����8�V����8��R�`���q�w�>I����:�4����i0�R�QD�����ih�s���?����K{�-I�i��,*�*`�&?�:�A�@2���Õ����г�*����R����:�m��<�;5I�`���-���v�ٸ�٤6"[�a���r
�r�{K���
�|���$0��0̩����6��G�Y=��m�|o�r�[�߲�]�v8C[�Z~:C�rL�I�$��������N�Ͱn@�Qks�~~S��J�):�a��e�0��?���� ۮ3D��4*V�Pę`@kz�����.N8~��#�jֆr�^�ˇ��
����z>��m$TԤد�b��z]3G���c~��&�t/hC�+E�^9�lk��P�j�Q���f��s#�X�;t�u�(��H$�(z�����0.�w���!��s�%����)jQ����;�N�o�a�ǉY��O�8f@���ݚCTMd�澂������~
fE��$~��h����@\j-<�Z�'7(��I�urqB��\����%�
�m�z�\�>G:�|`H����K�Y7��\?㦿{� �bJ�r�e������v$<�D0�LvR<�|��Ӓ�>�a�i �@@�;���&ղ�p�|"[㲙5cǵ��,G�$���^��^k�"]�_�YnSгU���|q����yL�#��yԁ������3()�"%c�.715��%�+X�b �)�(״�ڧ���`�i8J���}ٔ�eŁ�pwD����1 pp]����y��\�DK���4.p�=X�jo1�&���j� �Ab[����4�٭N1j����K�9~L~�Q;�*X������TΙ���F��7���[V7 Y�꼾On!iZ�jW��x`V���\�/"��\vo^x��㹷BG�����@�LG��=��X�0�. g��d�] ��/n�]s�A�P��	0yt���WGNJ^B��MՑCs�M>#���Ê��?��JG&^�A����wУ���p#@�-�e��A"��W4�`v��J)�ϑ3z�R��*v��8D�����nB���s���d���̆�<pҩKB���̦e�� �?���D�u;�О.#�Z?Ȭ@v���p����F��lMm�0�>�]LGs��'���Fܸ7N��{؅nQ�W��G��H*�U�ؑR,��P���T�B�?�;	��[xC��?ؑ��U)J���'L�yў�[�ز<MQT頑�Pn�԰�3;�%��#���,2�#�d0�=t���ZL`��M;�B҅F�b�o�_�
7t5_M�-$0�s�8Jn�!��a��G$;�@Zw�.a�O�����b�u���h	T*	A�!���F/�F�X���g�%����VW���N�M����x��J:wrz������Y;5.�q?���V��(��,��_�_�r����ѧ+tq̡�" �m��6$K�<ɞ�x��x�@��UC"�4=��h��������D�[Q���`�q� �G��@<ܼ��Z�1�O�����A_�y�θ��G����!/�1�՝�0ϕ�ӕ�ߊ�&a��L�id�W�����L�c?��v@�lC-cݷ��}2H���c����Sq��o�s{<��I�5��H}�
��WNo;QN�0g�v1GN"��h��,������m��|RIk��2/�60^���-:?�5�i�����?�]�P`�e`P)�J��TPw9lh.����풓3��!��{�0z�����ZƜ�`�mr��ڏ�Ȑ	�+ϗ��������^Π�&ۀp��R�=�̂>���i��ٸ�� }o!���J�yl�����~�hֶ��x��;PK� ;ށ�����n:����4�~5�d�9�81�{��p3�FX 1�}���.�y�������,�Mp\�M��ÍjaN�;���d�9�IWj.��x�3Ý��D�A��'�������u�J���$���!����ݓ��h�Η�i{~�Aç=�/��w�iA��br����rj�ST�1�}����q��Y��ȿ;Y�=�7�UE��XF-M�Y*�mˠ��������Q��\����,�"�T58�P(V�x�R���/�H#,��f#�e�rTxX
�x������L�䮉]{�Wa���Z*r[�s��t݁e����첲�!P{���[V�I��6d�42��M�k	�_��u�x��#�����1,��(˙G�� �c[]:�㾺�Q�v���ZR�{�țuK+��G�� ��^�MLK~�OD��B��`)�̸=�a_�+FqtLj�\K�3i&�K���8��S b��⡽'�$k<0B�J����4��y��s0@<'N��<��.�8��{�*2̂��9;~UA΂�*sTc�L>�mC	9!��;�b劅;ϖ6��<��K��)e����d���K۲-6�#6l��ds��;�&�49�\٧����0j���ر1�#ԉ?9;�0�0�6qP|\��yp&]����:�}�(ɰ$��g�ԅ)͹@k�`�Bյ6�S�������5�u�?�>��/���I���o2J�u_�Z����0����r�4����f�*����4f��n|�7���{Q����<%g�#�35>�_\�m�h9��+K�~� ����/��f���+شq��$i\�P�+�e�~��1�xˡ����B/�b�n<���:"�m7����ʗ����Ð���b��((����
^4�3'Cb�Z�(�׀-� ;e(�{��
�Ț�)��)��Po&X�w^����Q�����$[���]3qK��E-� �H��Ë���\�Ik&�ㅒ��Fc��
�|�qLY!R̎�=t:� �9�3��ٯ��5\N]��
T,H7$h`޼�F�˾�����d.W2&��$ ]��x�WyV%窴�/ﲼ���m����._>�e+/r�ܴ�u��|I
��b`�':7�a�Bc��TyE��%k�%`L��-�f-���  a
!ZY�*���b.��Devl�|��'6??�?��������C���/O1�x0�,k	51���c]��N���/W1N��,6��HX�>���~���������Q�],�j��v!�iǦ�\��4:�+&��P��[?{��ϓt�m����.f��Ü��2��٬)�|n�-��q�s������pc�����P�"rt@ ��/��t;�ps?�	Z��C�1E��ӫ���Khe��*u_����@l�V�3�%�;�@dD���_j��ˌ`1���J�����0����/�0X� >���:=��1�0�;�=�dLj��
Ht��K������9Xci�0��V��VV�v����d�� �vQԀ��Ԍʣ���j��8=�!�M��{��l+�?{\f�<�N���'���#*%1�N�#��e����2E�60(�E7�OR��B����\UL�d9I)�]���ew�;��W\A�l��&��rcN"y8�{�w@Z�Y��d�䖋ŉ��;�55�8]���U���L�g��a?F��vj0SU����i��LCTf��t�@ٛ�㍠�Z����4w��,��*�m���X_T⋏����󂭛i J�=�K��tf��*giƂ�q�EE/�@.~	FqI$�5�#�;����!��NL@�$�19�
��@�⊡N%�(�H���֏��c�P��#H	R���Jl�H��S.��� ��BKZćYcm��q�̋ �SnΉϽ!�x3��"�����(\���+�x[��5�`x�|�����*�����^(��A��9b�D%fYv�L�iv�%#9�O.�ӹW��L�rq��U!�E;7�l|�fV�7+�.��Nq��-�_��9���#����{��8:�O��/Z漏�5a]Y\�����9�~ N*e|Ԅy���:>��~�M���}q����T
���l&�"l�t^��ִ\��j�.�[�8��S�7F����·�����X��Q�n�ݼST򭑼:h:��^�݄���,��a3k���_�\`/��C���
a�i��y@jWk%9{���2Q����Qh���ynQfa���Vf�ݫ�"O��@u��i$� �ua�B�A�Lc�&Sl7$	L��Z�	���?f`�O�E�vЏí�i@���\_���mE^:�(�յ*�_k*mLno�FlNR�,y���Xw!W����N1�G�� �c�i�6<���}��o)VnO�W�I`h�jL���BܤB;�
��:K�}}y���TV�m���w$.D+�t+�	Q�����i"�V����ӳL����#@�~v5��?�r�+G^�7���z3�2�h7�r��<[�&��������I�ԐӴ���dSi��q�*�W�Eio���Zρ41�bIG��.2�L�����F5�剕B��C*���#���>�(����Z |��^o�1�a�Q(P��M���qLIU=H[<�6��(�&P�[��;u��P6nf��pi�Hǐ[�yJpp������ g�'*�k�¯��.@�����+�n��2��R�a�l���2׺�"X��w�?�j���J}�ɜ�#>�n����ha �h������)@�bV�-%"jj|�0�G�±ĝ���Mb�����	��k��ü�c1'!w�UZdď�o��L���f �%?����! ����_G�
y�(���Hwoԉl���߇����`j~x��.����?������K�җ��h�W��(*ϔ$�ݔt��:����Uj�.��ίW¬&��)�%�IK^"EN������R$���ai�Ok���$�M��?����>�x�J�>�_WL�ԍ֫,Q@SZ�Ќ��ۛb�i�r����u�������=��,��?w�mL�,�7����\�\K���}S~z}��������Ȣ�}D�R�8��<��� �y��±���^��M�p����e���/=��[>�Y�_�M��ӿo��<��%