��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H������N݆��Ȗ�����}������XQ�ǔȀ�wu1eH��F �O���6���5ig�a%���5�Ќ6\�f����^ŶG\{���6��5	��p��S}��jO�@m]�;�ˬzgv��4�i"�d-Ψ�C��2�g�˰i����xW�2���g�~�E<�?Up��%����
���'඼h�{��3�ThE_pסsKVJ�`�jѺ$�x�5��-َX)D�/8q�]?�|�b�GS�|U��#�J{D�|�?7�!4�gUnK�(a�5[�YK�u�|k���Z�MI�6��$�~{˴�B�Y�K%ؔ��^�]?�tڑ G(v����=a>pY��������Ԑv��MK�$���mhy`�6�d&�{ќ9QA����*���#w�@d�d��7;�/�7|�E�i^��5'3�I4��u�i�[���\�!ƻj`ﴱ��ޅ�/ �IWƝ]�]�f3/�B��c��WX��#o��$H��SٗK~����C�,=Ԑ���N0ћ6.��:��z�?	#Wv���<Ę�X���B�A�+�̚؀C�#���P���g����KT�1H�t�P�riE/��*P���).mL+�I���K���O���|����	��9�V�"&Аx�K��)�MK�J�l�o�JE�������Y����Z��[��E�\�܄w��U<~d�~0z��=I��E�j��J�"���Q�-�L
��4_܏�-]��̖ ���(�� ����۴ ���:�T3,�]Ѻ��a[ �]�-p/�	gV�Xa�{<�Y��jo7Z��'/�������R�Q�XY�(،���U��p�|���f}8G�6��O��\�(;}�[gy�����A�x�8�-��w����K�ΔQ��'$� �ߑ��9���0�߻m, n�P��&�ۭ��:&f�m�}|�O���$�USK,���u~����i��l"�� +��T��H���	Qx�e���YǷ>���jjE��br 7%�o��H��%֬;Ci*�Se,{'��}���p�C�F��y��IT����3Sx2VP s���V��+�"4�E�;��5P8���Pq5�Ǵ�1����I�'��2�+��ɳ��{'���y�����]���a�3�6�&�0T����.J�qiA�w��<�Ñ��fy6n]���^FA����4�yKm�Jwdu�E�@�
B*sF=���;T���Q����M�:Xe2�D��Ma��\8I]t�(�7���?5�
ǀ8�ӓE.N: �˛e�Z��O�\чR5:^��%Oy}r^R�bT�eJ�&D���> '�\�'�p�;�'�m���R����VY����ZK$�DU����˅���T������O �[�ch���ԛ�̈�����>#�5���e(�MW���pc��9����s �����il�Y�0�vg�����ղ�"�g�g^Bx0�h	�,�d�z@��4��!i�lr��Lm�/���˰U���KaZ	!�1V��d��ro
j6�Ivk���.�ɽWU���Ab�ŗy��\&~�o^�g�di�v�%Ơ�=(Q8�Ra��JF�$7��,�9]�la��oT�^��g
��R}��ot�.�=-�p?x{�j�N��L�'E5z������̯���VY���z�!ed�_E�I��f� 
��;���r�qmD���dpz�
�$\v���4���z��#����O�(���� $��E�{s��UX}�_9g_���G���ŕ·����	��M�.ǉ F�ji����kU�
�]���b�I;��}>����X|�o(�e�R��P%r(�Q$�Ot�AU@��nt$6��e�n�����,f'��}r 'ш� o&�p}�VT�<n\Eb�
M2��rji�_��o���7��H?��O!t�M'��oJ�*���)Sj�B�sr(�/(IԘǼ?eO=쀰�g�&	�D�����Cy\r�Z�@Ȯ�:��LT拓Z�܊m��Aq{u���䔵|R�����!L�#��)���y�z�3��ߗz6x�}���F@�}�+D�H�:R�T�����������ڈ�d?���ӏ�TO[`X����ѝ�?ѽ�ۣ� �/��S������r*�r��=���5��ݠ��� X?�8��uW���-J+���F�>r=�o��ш��ri���^!���g��\E{�6Tth5��(�O")�Ξc�6_؝h}�M{��m���&,w��'��l��5�C���MP*���Q�)s���Y�:�e�5碛dd˘�3h�$9������S��o�ᯇje�{�'n[�E[�6��HI���SU��;���� j�) 套��l�$��bC1�%8����;G�3��1!��7�ܕ$3�෹d��Q��O������&�������X>�����v[s�26W-�gШ!2��&p(��yX�n8+!M	��'��<����&�j[e��tp�����dp�+Xdr�1���Y���D��62��K����5�WІ0��(�9�Ek���/�e~>�6��N�������2J�B0	hQ��T���r�E�s��~�ƢJ��k�؀%��B�̓��Cr�_M5v�*�[��S�
Ifn��.���d��ߊ�3=�IyQ� +w韗���LJ(F�0m-&�By�`=�mv��~8�0�����v�"�j�E͞,��	�`���s����'��	w�\u��s@�\c�u~7��'��A��A���z;�:T1_���h<2�ޓhM�v��&��!3l���Cr�$��\�(����M��ә�>(��BE0��zAip���UpZR�*�Xq�v���j� e�v�����
n'�����N [K�6U�|�_�Z�e�}�<ivC��%���	"`F�+E�>�l'p�Pm/cଈ��3�'�N�I,�h3�3��Ǹݡ�"mHwڊ[b���<���M�̈\E��n>%*�K\6���3d�hR��ǌ�ѝ*u9��J�|ѐ�
GW�\�����7P�����8)Q��Oa�l�^Z#��꛶T���S��*�=:'N�}���']$�C)��	[��/~��FA� "��2�l�q�0���E��l	���Yf�.2_B[؈ܥ�t���3�,����x��T�z��e�B���x��T%���DѲD*�&��R���X�q��.��o~�]%
E>	x�`���R��'�`�z��MM}�o�e��ą��&�|-���H��:bz��[�*��E����2C�����Ds��q῱�p�ջ��A1V�.H�(��5�ŕ�Z�K��R�����X�l�� �#o�uop��]\{T!\W�с�s���E�����B~qB��o��l���Qb)����Ȥ�q���_%u��`�q���sn5��Q�Z���0?E��T_@s؀�`Kp���H�'Y^�a��U*�Ӟ&
^�̊��c!�gx�%�C��u��3c��j���ɯ0ρ} ���%K�>�����s��B���y[�%����H�g������"{]ÄЉ� ���.I�h�~4��]���Y�Œ����&$	���B51U��U�،gn$�C֕����aʪ�G��~����;G�*L���|?�ZhKߦqWw���Ҏ.gj⼑�l�J������D|���Q`E����7�Ḅg�l5� #��
;��&w�,
����b�NW�8��V��!L��nm5Q��z
�f����9~٫z=�=�bW;+}aE�� �=yф���S�q��Z4P�b�V���ך�&p9���>j�ܯD��#ׂh�0��-Oc9��+H��L�4y���!�mPf8�<�y
12�]��ο��é�cA\O�����k���E�S
Z�xQL?Y�S���S-�Y��k9�i�࠰�j��8��