-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HyEx85cUtoAuudSbbBxFNSxkB7g94EDV8hwQwmVvLLHKVzD2wRiduuzTScCm2urJl5AOdq21tMZU
QWGOVpZBav4derQLaezbW8vDl0iRkqBC+BTdR1QFx+9OSErD8Sd0TH7Xxm5dAml5dfVNmv+NQABy
aP5oaSVmahbM0N/G/24bQnMrGGEje+XzJOe4izDzN5G2EoJjNeBUooXR4qnzUbNwXHiv4tbaeWIm
mL7PBJoI5El0HSKEOCQ7ZdxF7QJTsUP6WR8CZOfCYeyzjIzO8EMj3AAYqXr2Do49Y0m1IhJZY9TI
bJqAMDrzWkDmubmToiX0xgiBDkt6mwFGAJ1gjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
PDFR4yjlyj8qi4ZjIDv5iJEHle1/4XWDG/o06AtldIYPlp9IT3nMwb0Eu7lNHhEspA/1+EGmLcPi
xb5sPyHNPiCgIsEfkQaH6OL+SJG8xj4JMDShDIJTzneCVkOPN7QU1/3bxoB4kqhJ2/kNeSqxcZUl
kNnPw8HVB7TSpYd/gw1wiqRAUxMoezhe52AWEucIA9SSDBAmbMTX8JsZOlF9+aj0kZTEn8Ov2C+0
Pz7dQ9zvNNIanr7IANL10KOdeBHoz1v59KNpCKLikG28Oc2lYKs3/K7V8FU8BZXPL1u7Ui1IYlf0
cLSWJm2ZT2+rrdnW2Xc/RWipDaeI6LMhrxQLMNJgRXxdJVYrT5RzIH3/XRn7kz4xrZ3ezn+Wi/bQ
FcW+XBmfNMFrNN7UE8Ew7ElqlrV3yzzIDAhwPQOA+UeKg0a5eHgylB4V2l1sLUDvZKIMeh4EV+Ux
xEoQGLAd64NJ6Xd2T7TJE83RWoQzjKwomlO4lATtdcUPY/BCtqhuSg7wWTVy8zWqTDhRbi2i2AsD
XT/9a4/TDgBF4VwofQu26aMzRWTd90+O9xYvuz2CX7wezOTg1nrcDVAy2zMmDn6VUsZpLFoHFIVW
oOU8eOLd7pNVqAnq5ZDLtbhFp6f0UbEwRmI2JrryrAeXTflIkiO0GWctHaLQFXXY3FPmdOH7pkl0
MO2Ua6sHJ+Kp4iguTtD9hOMl9MXx8r3MiaaA3XAFDNmG9l8PQVsS/QnnEipnBmdVZousWs0sdPN2
nGqMWqfbtROSCVvQ3lVnkHp2U366jLYJxee81vuHL3vsM4naJpA7RGPk+Y7NNJYVU5RfsxXrtWdz
ySEa93ND+cTFQFs6zIbHTH9d0RAGpws3sbgDwZ+vZfxDIZQzWy1CRrp7qoeY2xzJvpFKww47xTMJ
Zb2v5GKh7cPIxU/q6n37XjzJ/Tytzw3nTtjl8ePnnqysdVZfXk3Ogl5e6ieFTCSbzkb5xBaMaGNL
kvfBQUiVhZlSHxjFeS7RyNWS7dN5HSMHopLTxUvoAKEPH2Cury+4QxIsVK5BZE5yn44wApl5Pdwf
0eghT6dNVKR+wXWGOmLY1UstR39wHM16lp5q1QdXjT9VhMqUytwctC99M08jrL+2VR8Qo/EkLIw6
IZF2RU2d7nBctBZUmwncvLUHSJRCwcURHrIfJ6YgqULIS2s7BYvA2hghXN+sSEy733LbyiU9rfGc
t5AYJqP+rGIIqRukT078TG+tDs5BI/cRhwcASwfKVupbm1iPs3J9dA/1d4IKNm0o/gwV5HnAD1TN
jUBlSJl8gKI8sW2C6hlNun6zoWe/PbomgWYU8NW2xLgEk8ECstRyq2ax47Qzcj0kaFZSY1aTbkyS
0bGY96oDvax8jP1Pr1YI9cemYUOWiStDCNeK25Z3jP7AdOxqnI9kOY12bCZnDVQH36NLKyVap0rc
j9XhtfGDzXg+vq+/o8cpdZcVpuWxlPtQvdt3/yeta4q5MbExV/kn9ai+uchGmWCbXCYmIpjVPC/E
6VKpWq80Zi4AQRjRU9fXGFR04h+asoIE2uVLgWaRWz0/Y0B9pb2HflOB2lkk0o1o3H2lCPd8lKFt
XF3xEMwuzCogKWWAzBwu7JzMWXTCgbeQr75B5u/RBnFDpsOY0URsjNRoXhW5+CWnGubxcSM+Cp0u
jBSLbJSXZHAb5gERGHmLfNP2Zc+bbDWoLzlT26NqxN4ZXk7yDiBFFdFLUXeMsVmvSdbhoZerWRdr
Ei/qRn1CkjKgyr42uwBI6P/h2IRFxnuIAAvqwMh/xqVQQRIQQauZeGZRazR86y8Oqj6dmvLj91f3
rPfqL1Iqkvw5Q3r4PVJCZ33iVkh++b1bvvcQOXeWUj9ZT66u4O4AhrKxUPoECK30qN9tviyqylKT
iXys/U0dGzUaNDKPXQmwI5LDSb2PV3GhdS4cmXP/kOx1kb+2fZd+5OXTXVwLDEWtgeZY5ih/yn++
iz50LRyI4hKHIL96vLfbYpY242Qv/vsa5h6AbqFjFBueY82ZbAxzwag3U+rGZGUB+JcM4/CStzCW
RJvB0cyopa1OoWGHufFjYs/qQtOvCwW0HhvxZLDKUsSktqUVbhbZJCW2+4f0fwa8R+YL0jDwsskB
3AkFfu+Nr19u8c77lMTPchcsgh8jJiSaBNu8X4alR0nIWgEra9sCvDQD1tyYg6UQsh3A5IgBj91M
MYT5RZ1pWH1RCij9/3oyhfDXJ5fi2sxHmgIttlKsiKJEScGcgfUgqDE0oXEYdJOeuKSvzXwyaHAS
cjkXy+dssVh8jc2uZcwFJ6a21VLfv/d6BRk2Z8MJGMF1KFY27NPg4UXSK/wyGQQsR7TJwcCcV1+g
ZPFlSc9hKTzv4AL3mypFDxxblhtl4c7Ca1rc9yUDmMbI19R7fxOgGAKjxRxovbqFTONqlCvMDbqL
gPZKuOlE3MvNWVhiTiXf+FBuWVdVbfHKXrE2S0rhj5ZZsH6cd/bt2GIFzasVVJrab/1ybKdkHWMN
dFHLZb6wRTuqVHTHMnzkV1AKZsvMbeyp9u7fzEJ7hx0BuVTKUUrVdLk8YYqzivBmm2fGrYvRSd8p
06IUdymjgIZPkcZo6zXWv0o6bcCs602gAMcsiSRGkaOh2Z4cgcXI38NFYiEJkAkne4Qf0oPMvl7Q
XMUF+54dlJlAiprpEfcvFofjOMGStywJKiOAVYoP3eQklsdo+UvlO1tgbCdQgU0tgLKW/PdBKIS5
qQ7yqm0AVjlUL608gmaeGawd3ex9zsk5+HG502kPBFkfFutZSAXFpkntm/vkTyH1nVJxv+jGL4K7
SGBI2oNswIye2lTD+pwWYcdnk7oHOw0EJn+Am0QbsIbJ24AC35WdSycIYzbCRgjnCiTZcCS1l+VO
pBPlWCy9K7tekqPzHBoCroytTbcjAQJ7GGxWSOSMEeFCQKFWLOXETe7LQ1zGNEf1pE37YumizoQZ
zvGMk22pDKhJGaHvLFDy7QBrIrnVw3nNRo+E9fsMifFWVzwDYFypNTJaUlFHLKRjrTR0+xKCoeMG
cvUCHBN6VqVO2pJ7J/jeeWKg35RmoMVh+qzmI4puFnOq6cqf7n/CCNfWk5QhUGx9Ox9y8x5tm2KL
N/eCO60KwXlaecj7HfC/ALGKEUmCvPdlhHBoljjGP/Wx/0CCPZqSv25GSrolwtHxW4ACd6d1f3On
c2wVP9HD0iz/MsQG83EjnZFGjedy1HtVia9dVkuelcTfYqIk8M5lJ7lnvPYeiKdsSXuSPQNIvWcH
hQUJ37zOprLXec7aUZlrR6CWmLS7wHG+gZQjlKoXQafP2NmIPlmHWkda187LAMy//IeSV/vW/PnE
BoBlB2D1sjv08RHVu7GK4KlTKM80uoDhayLsjzgwBk4KRSJNtk8KMiz1Nr21DSyGylbBKNFPTndm
olseAyzOpYWSOjAlyv34IeHCbsk8B4iV4KFZjtHMvNLQ/BBRntwGboHGHDY7kv75QZt1m4CH4Jvb
gvXPhq56/Gufc00D3iGq2jIqLVEOM85Yl+dmeiUvzbH10iJsfmFPshDvOx6x38CcqNlUiYMtu+kf
zc1utW5Q9IGgi2gBBxWu3G3hTA7X1t+C3dyPc71EifttLlN8gTLfQXp/J1z/4Iyb+ufs0YG/axRJ
EOYs07Bk99AqPzBsDNNQu3EjKLp5YD+HFvRzVX0stZhN7vEiMI7DuMqoy5kewYea5EK4j2JnzvPI
6vMXZIWfEjWp6uCI34k91vbmRCyUXCfMDEXHnyLkBbjZ4FNMIFkPGPu5lYqF3g0+RwIw7ObdnfAi
rPpzYBZgAwAk6clODmk+A0/uKfqsvWGba8iEKVQzk3I85Dfu26R54tIenjTyFF9anANjH5BeOtyP
qFZDuE4+u0lIPowlXeILbIXua+N9InHv8aEO7/yC2+JgaMRB8MkhKfviUhHlZi9w6Afh34gEedfY
94CC430EGjq4yZB/Y/KI+kYUQL7oMER1yuB6NiY1POcb1nVgmKGt0R6LQEohJRcVjm46iE+LEjnL
Es9RZUrJnzXjRjQJjhf6zBGQd22y4Ylr761NOnZQP85YolPCfv1eunEXM8zB5QlwrYwzRVwNmRzt
0hO/eEdUE5VJk3uCW3RRe71Cq5I3+GGn/KJqCAsLUoAMZxKucnId2DIKGef0lp63QYuyfUfey2DG
x0/C85vgcQXmQRYbC12cfttkJvHFeqy2u8IqC2FekYf7wT6TVBe5sLokr1c3BY07a4O+iqGHLWP/
eYIY219beSdGujYba28P4c4lXjTBaW9yXM0s1PpFkews72NrWVQynpwzWStLu0roBT1DGnvWYhLy
1dQ3+Xb8vDTdOldqJBPYWURZ3K0UZXpRKUNihJKZVX5LyUYtuRZndYshCpNnHQBLl1KcQLa8HADl
WhHn8fbiPNrwZikZenNfmpdgCsOedV3yTa4aIsSluo+KWbuhQxNCI829yShqNNf4LEPI8OMQsZeO
ecpyEnj95K8m6/jgUbHLQK6Li0KqZTJ9h+clNcXp0h8PxjkkZKPnakHjj+ovjKWziHEgCsGIe7kJ
pER5GsHWRi7aE+kqOG4qDgtBUYZUaZeBs97tr5J5llfCPv4ta0v8wKgTP9tYnPEN9SdJtvnTHdy/
kl/xZv/g6Y7KkHweEz9m64i+95TKrihvdqj+q5HQ+lwhZgj6Hwy5JDfgOOCAci5Jp+bhcjTA337N
r2oYTHSDgZk8ZEVfKQyDtWRhvvLYYG9Rl4guyheA1QQjO6ai1EULZcQhtoIownx8d0tL7oZnyB0v
UN2+BmztoIUvwjOaHU2oRE+/jpipiWoeeg6mWiN+TZLCHT1Ref+QDP/h6eGy7FI0Qo/Os11yGNGR
uOBIYex/tZRvYOnCFolmQmrrPNJOo+zzfOL0EvvvLL8fsj4VA9S70mTqo7TscGbt9kFbAk9yjBct
1FfDRFfMdlpGTC4700bc1x2AP9JSDrGGHxpjE/liRarn+I9x2kU4nOy3eLiyObsNx2KOUA8/8qOs
TPpkKyVl0ZQAUqkhcxL4J6QbL2LLk+ZJxCYfLyPyjgdo6xNLgVLjKOpFPMPG0iB4tiEj+QK3GiGn
9wHLrBzzvzhX20H+R+CJnyH/XIptLSJJSNLIHMMK7kUH6RqqqyPSlWXW2sFoSuMxsAU26iionpCw
s752ctjPqDwOCvsWHfiKh9kBaC38ma5+qjzd7MI6PLR93XhsYZFJoRZoDSXwC89RJkc1TeHuxh5z
2baxco486OSd5QlBMh3S2S0FRTys311TSrM9066FAQy26fqYSUeAQHagdYDNyJcjy5ZachBXnYdd
obHcJwyi9kAgzRkHwWk3S62KNLasXhlsgmp/jb23XLsyhLkYWLJZq+KWnYi7cgqaqE4SPKmh4jXW
E4QfpOM+EhbLVGLRYIFC8MkSDRrYNfWSB1N4tUSz66ivaBr76mc7ogoGqxm0jh+Q6dU8/S3hj6RI
Vekon8dsMCD7yn4UKBTpvf5hHov/d3G1QpAoBsF6YX93kQyZzDUkvy94SOLUf21G4b9/BRvDt+K+
HoJu6QEMrfPQzvSQiytQsGWgdvDdhNMRwUt0MUuIpEMPKF0G1qbk0BobSkvLhW/tgk+f/hg368Ie
7aMyPgZma1ipgJNVL+DTpcm56IYNggWMlUr/8LQ27vWlJXXLiNxXYuskGe2mOZcKLBzoBD6ie3hr
2Dl0srIBIwqZKDDMzza35XlUboMK7tG/jEQnZ1equX3wjjEBSMaO2GaA6gRE9phKzuYZM65vm1YM
Xy9OtI+ock8V1alKF8Nb0K08MNpp2JdAcZKbkfKSuGyYfRYsbrcopKLbmR4Q0OEAuqvcfpQq4rGk
XYxD4qfK6S6/PFkIwyErteg6Zl8c5czXaCVOeVRYBAqh4mwERnMRgSj7vMMOmyCfRW8iZjWfvzu+
QUOSoGDk+TwShG8Eoy79Y10U/trZBsRHv1w8+r8nImTE3jXAo2qu2DlE3pkqJyaCtnAVRA4shUex
x5p0jxZAmDo2P2s20kWKs/8jhs+FJh+Q71wJqHXjrHL8YFqFM63/sunuVKKiOsuWgIjDWH9J5Rmm
S6/9A83OEwrsqFF0La3o3OM83RJfCcqRVzQIFi56BKio9MWfY0L/zrPl9bHWat5BICdGK/kmPtqd
ODQ3T+cfoOvjkelJ4N55VRv3bF2draYBuaKXUm4Ky5+xxvZokGKPchpnci2S/iwgznG7U4JBUYkX
wLnq4+B0dsBDvG7YQ0LLabIK5QqlgWejpr3AU1hFrJUss5EwGlb6rjKWRBiVAB/sca2sjUZ8J+AS
VoFyPB7TCTd6v4POJ5dcTWpLq6CMtAYxuOd9fT1u38tpQyzQB2o9aZg4j+uO5bE3ku2t0urksHaf
FgubY9T2j00TT2Gg+b7lT6cKhDLVqwCMpLKgQqTvdzhBN/5BBSST5VwsjL4O0s8oEJeDM00+ION5
qyZ1yVChlsnDfjVV2GTqAVNVRF58r65yty7JkxkKwl7ylVZy7nLgH+su0w21ACJ+24rkw2pBIsrI
5L43YGhnY8NX/YYgHv6JztnBwDPmINkSadVd/7a35M/KEQnPWsUEL7O4hrDR5v4pCEUf96w911LW
HxmiSaiibQrgI1cIB3Pnc2wdCYXCN7ACBwOzc/rlOprmlecfMZwv88pG/ya2Jl0rMHVoxscIAOXJ
EI6U7rgNtnFKbHFo6/lyV/oBz3I6xBsJ27XXDhJjfBXVBFashS50RJMKPnacBTUAV4TlO8p+cPxR
NYqVtSXX1fYvjXIYQyF0Vult2NYcSEWQQaWuOb7FJrg1HiFw43qbXWsxcyVyigaqIZ4hen4uE40K
hRSVUaEOMHnloAYbXMeK2SWQi1Uq2/TMpBHLx4drhgTknVUr/iGjj0O+ke0pn/F2uExuqR8DlLKj
peW0dnxnN7D6auPHedCMpl4Te+4/hVHL7MxI2LoGbIThrHiiT4x48pTeKrUGtU4wvB87hfOYlDK/
oBGNL8Web7I5BdJzRGRLHhyuv1HQZAsANRl71YqyF0UUeYxksNHJlvE++rO9b2yeJTr/tygZstZO
3k9TgbK5HEfuRnrHfdkDKllczLeQ4kiMoJk7Z6TZGv1NjZVpz9W+uzklag9RbDjFMGZPzwCjaMRJ
laRFfIfdY848YXKUCVJnm05v0fIFb4VjumwHyEgDDdOmiM+CsC6HFLoEB5FVyhBBiDUQ85PpBeir
cC5TBxRKkoSKRFw0zmhdgmJszgU+XvYmycwFE9YCo++Dbt5t8K3AivUX2OQ/YnEqfFpf3b4S3ZPR
5Km6Zq2Pj35dMvoTqQqo+ACLYjWD38LPojp3Elrsfn82XuN0q2wtdLxGsEQMAofSsMMaE/3uCUtJ
5frTaQVR1XPlS30Cide4RfzKAJQuGOjQxspIPIS9p9fRc4dz/s6fmQoo1qrstI8IKsOE5AfmPS2k
E67WFrKVhruIRdAZwKWqps1VhAGePODp/lwM8wt95R/NV9WkjS7zt92II07hvYRkDMOYsl6kt4L8
gH7lY7abLAXuLRHCVzui1vM+BFOyhRxeeJeHAEiK5f7DbsogxgyXYmTvN2G+ewFd7gJJwj21Qx7G
RkvdYpzd7pb1b4ZXhUpcgGNM4/Lw2tLZvOVHlOEYseTzT2wOCHAa4enXNZV2/UsaZxtIGNNeFvd/
G3WB9i8Q5nXT+HOJixb0BWDVG39rucjYULg3toHI9VN+1qJD4TJPsgMqS0lsNQYZN9MD+R8RxT0S
5DG86eEP77PvDpn7AVtxKJP3XVWx6ny90C1hghUxJB4tggZL88xB8nm+Ur0OiNBdZohLbfPZWfFf
WOcYQMazUw3WQEA9VYy3HrVGuStc3k4dCSg1RBZiswdSKVyRClr/6SRwpODPN15YK1QxVx//xljx
AfOxT1ZHeUpQCp3107mUSm3N4E3x9386lckolW7qKYV9xj0jiziTRnyAGNgknIHNrfZ8Et4MNtAK
M+R2K1NhG4mo/hWtT1ro9nK1KNFzMt0OeXRF76VImVJxBFfnqs7aGPWoun7jmenCpJt/fx1o8yhi
yz2exhJtQzwRLn0eL6JJ07Vyk6R07GBg6u9xsrOIUa/NlYtsI6YGgWrIi37nz4/0c5c4+q3i1k19
1MzH4agarwkBzg8fCaHlsqoyOB3XvxiRggNKpDcHH4h08MhuyEbrBlDgjrDhd/0N/bFlHZZGYIif
hxdXXttDhXePzEoFMWrmiuWbNPsXEIDnwXfu7Q9jeqlTzeYORZvmQ3mU+aYiKo882TIuvExmvC2O
JPWKZv5k0V6L83pzABM8kamZrboQB5rwFV+VJxPZRZtsby7LDNPmFblDt1Z8HCh+u9mMmdgOjG35
kyB1ZvpXV8h1i9FtGpx1QZ+WbhLccVcQUwuaeVzCkrucGKuE+uEUgDnscizHi/zA5YyKVkAl+rzC
LMyc2ziAs4SEE7CAB9aqMn8CkpOwkwdMYDIYchMKmhFU4Xnu6IBd1Tp4AW0BjVea0E0VGu+1A3m8
YESJxK1p3AgIDBhc8IJOJynO2PIVHGLNuBVYd232SkrOs8Ad+tdaxtWDcmypu3m2HWnoq387p0JD
VYQdvLEppHNCEWiRG7pUgO9Y/rOZwXcRtZkCurBHhI3n5rSA8KK09qML3dwMc+9c9ekDs1AahpFs
mv5hZ0WJ3uzMzvKYz1xUD7oNejN88MHFyfauCUuq0gc6ENnl3EZangrDy/TNS84z8wNkKCUAeGU/
+0pCod9SYw1jDbMfcu300jhDQ5qW75GhEZIcuRLIo+X+tdtLXK59fzkm/Dvpgc9QhOOKm9W40Psw
EvS+sFUSca72JdDjH/YNkIGVGfm+7vcSZY7CRFimK+p2IVdrBxnRCyGkJW85b7Ik7T1TlcVVSFjz
Qogx6YmTsdmDPl/ZBzAyWPKEsVufPc6Wt6V/4pXJA6oy4Rg7E6/F8tOI/kpD5nYv518wkTtHpP0r
odMurs3bG9d4+2ESrZKMdhFtKnYn37GJKFEFENTD5sOqDTAJb7hmexqjaQyhfh2FBaytJ4NuPO4N
XGOsiV63UyWzlqHQxy0uzX5q4Aq82mi5a3Rx0Z7nrbKjHdZY9BqGHYYyeEZJopBbfqiVJrz0Q/g+
Qn7o6Lix7MLvxVywbWdOsd/xPQh3S077jZK8h202LQyFKmOatV0PWNVxqd+s+mtZ7pZk3WckCYKk
CV+FfnxEwPqN3nt0QQF1Ur84KGbhi//mqauBok4zEi8E8N+ruBetfb6aHOS/Qv85FT5L3QQmBNiu
vGXmotZ9DcqIFFbtdcGfO/ctmXUo+Q+hd4yp4OHE+zp8D7ian79t+1n7TAXDMpOi6/DDup84PmhN
pYjtv5AwheXVW8smUj8IikmNEt7R7/C4oqRdmYqacw12dVNuZiN5ECO2qvfc/U9k/nr2r0elmpba
yR2272nZzlys8pEWuODVIoV/nCDFGWrgUT/BxNxiHI351DQpQya6naA4riLlqymThzfgIsBnWiW1
LPcVLwKOr0CFgPCq5406vtjqK/dNylxA9lT3rwtcUEaTH9ULPOmaoV/T0UmQaYqivkuOrbN4JJ1l
PO4S3fHEzRMfmByQU/3695AXGCl2H1+KWmXzPEGstyNao4lRDMKotU5OxroDpirNRXXi5Hi8ZcFB
7snWDTsz7nezzSB/E01r3OsuhlHXuCdEmR7WbZMHRgNJf4Lfi8gR1Dk8+ido705cZq2SLo8So02H
oFhmSTK99CV5t2nUk7KFrQsu4FxHLwnJ+OxfU+iPm3yWD6sbyrLGdO7m1sqZAuJb6SGDTv1DxIXl
RX5r4TNE0f8n5Nf6ihjWLwKEPyB1yFX6CwCrB+VddKrS5yO2EGARRXw7t6KbMKmsYViGMa6IzEyT
XYMS9g1Wi2dro6MlNUNbAKZmXwrz0PPZ5gFRIxvfMm9L08f2EbnwHaOjJd0tIo6tKDdH+WIFpZlU
4Xx0CQ1tlcLt/t/4bGgplvjtTxXUkPsG5FmwjezKBFQsSYt1VV8bcB/Rl9drk9B/s4bq8VUIf0uB
Do7zMrDiXts1qH7KVDlpn/4PtwjxoMJftnQuMxCA2ELkmIecZoL/fRpxfXXtoxSVnQ40n/+8QHL/
10v3FqjQuVO5xa6pVyhbVh26wfMbJp7bE5rTjSJaO7He4eAT9P2OAMC3J1jz6h4jrgBr6Ft+fkY5
W3/pM19FvMQCN/evATt87qq88gn9SUIl90f4HAE0IACWZ28G0nou2TQYthKZqeDcI7LCel2BewpQ
oRMJsZfTd72zVK9bM/0+ufaOw36rn6SxtWHklLE0Mzo9Etmw0miuEr+fPid9JGRgww+e9pfPwAxC
lSzXszIKgzw0cn8ovOieAODDE0/zE48EFR0kLeOckSswXyxO0slDNhZxrW1xCjBngFVVtglfeGr5
6z3g2wFhnX0X/3PuQGKeiqlmFTMuYYs8f3VIJ1bRm8lQ4xmml/At350cBLCLw94/zqB+OU4oV/pn
u/QEy140AfdNJbax/VjIiQ/es8d5Ldcd4oDtjFiBYNiiyHJBheuFSdBYsWdimNOeGCjiagH4iUfu
uC6OjoFV46yIOvhH1fLnqYPSzV42JFXMzPpQdOhk17HggO9mcYCoDCsFBy1sRly5aH1FFCPnEX95
MaJYVmZg9H1THy4kVfRO25P2u3kFyab/EoUoBLEshGVcRIW6Yju7rByIuFxAdrJNMgUYfQ/IfSPV
B6nFOAV/8HZxpU9mqrSFKiFBTrIME8ALhPOPUV3b/uYheyetsQNOmkzx21hDGvR0rGoJUX4ITBWF
BviLx7FqZwwJO3GlRzlI3hCc6rrX+OcVnZyvaM0wECoNFgapi1HayiktCgtmU0nCDN+664uU9Ehg
grzfmBH8HKIQEGdkHym8G74wnmooQ/FDGDHVby+IohHBmPOfc5+gLPVhrXBT6DTdiil05z2iQrDq
3EC0kPvtU42JRmca5g+b+yCDgyk+5XhtVOOYgu1KrwpKcN3WLDa8SzvIH5PN6lvhlAwCzF5p/K1U
kMGiqQSe8vfWW7DKRyXkEL2I6syT+FsqdPM8ljhKjJC03SEyWfQENFQyD3sz8HX/bH+Ta9Fk0b9b
tdovg2f6isbkQoLn5P59pVQAnb6SFOiiYBHVlYuLEbHBvq3EgYpQ8sWtQ0TiI3xrBLYiMksrmwVH
2EzWoXe9PbCMh29mdJx+phsFp18eEQmnX6iQ6CC5oNpw1Zk3kbCRIT66ivOogHkhnN5CtxpW3tFb
DI4O5zUsXUOPkiy/+N19bW+YblTLZoRG7UG03r3przRpPkqIYL9XnX6q4Qslj1VsoaEDbrv1z2vw
D8a8CuOWWvTHSWO+seRsm7s0k6PmTDN4K25bSAz9JybfFuFfTacW1FzQLkRDmzFpfSMhXmRx+CzE
0ycLdyZp6FahX55pGKtWmZAV6CUs/6gUmBvOJqVIPSz3y578m62uW/bnNJV01uwrApn4iZGBF/+1
X93NJv+5XE5UudtzdDP6DIyMtFPM/Po3agFpe1b3MUlZrfMC3yP9J0WhT3V3k/x9TYFPhLJPM8WJ
kg2g3roESKjoG2I9tQdG7W6aDBsR+aEIAAPwoX9av8hVpEGrlICMSzzSx2ocKLtyE0JLYPb7CBFe
YcjbqrjTKc9Un8/oDqr8bDFgjVeG6NOXFtbsDf4fwV7ZlGfBZEZaxIxwx49cbR0p+OJQGX3kUZMY
kj5jdNxNGMfzhbdupGcwFS1c4ztzQaSdIYjJo2FzH5ANAWMxaRUcZ/RPIg5oSxMcUekC8xih1pZC
xaBoy1sQhKsR4sPu3N/OBKV3ZBxSWswwfCKyHKkTB7RwatgwuB1I1erIU2yl8HAweoYs1G0asOgy
ltwWdB+wE2TRD2iAIAEcuemJOMAGfYKNN+JmWTHsVWHFxN3SH74rC7t/CyeaEX0LfD7fYtCWLIRz
IxxcD0uLDuwmB2gsHb11PAmfxY6+bxNjwf3bMlZ4kYk0Nk70Xx/3tWfyYxeZ9BE7kHcimKambHIv
xGTZw1tl6Ce21CLI3Jr5ATzCXlpXoufxL0zwn29SeMSIB5scT0hv4AAikcOq9ctD9SqSCHKPDn0z
RTV8OvpD7aYzhi+eda+YlwypEuugduxGA1JDa3Z4YX+gWgIK9Y/hjzrkQIJ+bKBghZNbjHZSl4zD
6sPndevIDXAswiboXD7EVjUVc9yX+btyWXYo0OB0Tr7MSJ57n5NE+P/K9EK1xY8FgWlEg/yfYjBl
lCMdU+sq8W/kWgyVwKBM+cqtBxiqMWo3Dmp9QSfusBchTx8XH5cE1xm/uu+HA2pPZtgQJmAStCyL
IPMsYbx80bouZkwodH8DkdNtjUCAt6+XyQY88j4PsNja94r5wdtw3er/tCJeaQp1VkUcS8Jx1J2e
NN7Gcm3Fzt2//JvTPCaxqMAfx9JpyMlTPYup/Cge6pho5Zof50tgoi8PDCdwx7EvTopQIGnxEcze
F87wuQRoeTZjEQ3EwqwvtxFvHQtRfqYVwSUZ3Z2lilQbBsI5V7mqSJGrSBVZSUPWYlMsVqAB4Lfs
hOmFwiGquSL0qi5QpYgSCvjokll/XuMUjnL9ojpGTRRsQatiNaRLYc7k8FCpPdGj3wPmg3AfskaR
HyzBVcD5EaO/WgyciDUSzEXuq2/WC7def8fShdphG598rTuxXTNGXmS6BOjuF9bn/cFZ05CfAlF2
SLhpYL6M8V7MDImpGynpsVM7vvq8nN5s73P8vLHeJ5TvynlLnDokxMcQElG+zCP+I+OJCqnmwEHO
LHtZ02xhUiLzXnbBCNlk44n2pnhJSLKn2KeZ/G0uofi/PI9yUhTAWfsDYnreWAfuaI5dt8EIn3hb
trU/vMdSCIZPtBZoZhbmlGD1sHvG/Nnpz9E++DBiBR26hD8wtmVPGbGVgAjoRQEGyXnoTjxAA5lK
EUw7iIc/24vdkrlaJ0L9NxrtB7u5n9xEREKyXWJKhVh9knjTHqLp8UuFO4abE6y3OKEat/5A76kE
Wb48SgyCfNhygu/Vbhbs1ZxQYzPMl40QVsHSX5XcbZXU6nATwUbS2QOLJTC7pD9f6IbYUOJy8xjv
EDsbDcT24n7o9y/jm75o7TaiV9CaOa+pF1Xewb/F38hQunihcrChQlSLC2uKWO/Sh3b2aC9NeMKv
cF/tlzcXPeYDSDIkfsZQ7vAfsT49a35qJdRxxxy5MXJwCSq7TQFgF1B29GAXGhwUSi5ozJfLXnpb
FkHv2sUDlTM4Qec3ql3BNDnQrNjVPnzWt+d1U6C/AXALW+vSzmbR3KP/c95Vjl5muU96Zu3mGzF+
iwSnfGqzh7DCmRuN61fcB4La0uoeaod7npq1EX8xIRl0akoIvwmakhIBDMZOP3IXqCbeLTilI+9Q
DMDXH3oJBKolUy41Xni3QucOEdBjQ3JPvNSPqTQ93QAOMuQz0f26oIX6tANHkQZM9kju9WSI7VGv
dKC7eK45/iPTBKMYLvRPLrpOuqusJdkkdtRs9d8E1i/rieLA3vbIzKxS4FGzzNWK+CkGU1Rh073y
k8GG83HJ7FDQHWeii8ZQY+gZDKYJyGT6JsxNTWIKYnn95z/hMBzJ2tKNPPydAVprqWxh7uO5qT4/
5T1pIUxFqnkDEQ4uwUOsbGmwT+g98W/vBIDnBhsuZnYnkcwxj6Jv6haL+0mnzCsLOxXnxurap/cW
A7ld65b/ZgcJOoJNoCS2p2J2HqMWXZ6Ti7iOHFtICW16SKmbz+fDrj57jf9eo3nU9IcjwvY6sqKG
gzm+nrsnfoqNxN6F04PQrXReI8yaCjFRLP9g75NEULsCXezvV/cQKQMZhg7zUJtsw83ph98zi6Ls
LC9kiOTcotArJQESiYdFpfyj2BzXoeZNA2mip3nmhdRaoe3mFm7lAv2gmSSFIilaqS8sOFL2gG+5
BSYcYho+m4rPM3X1ruFHfkFCZdd/zZFptLkHDH2aadgkG2jblJ3aF81FAHOkZwKao8S14Pi/7VRw
eivIvBUo+C2AqoFROR15I4GBHMsnFq2tf1ADmp3QxuQGQrsWe7ZBNS2Q5Qys3fyehj7wVLKyUFQD
l5gyA3qwseKm8zhENLLkab0yihBrg75j2uA1QUMeJNTsHDTYwxMO3h3schOodl+acEBjDYFU8K4P
tgztW7ASbNb3qM9O1IAxVnkUxcDJ6KWPfGzv7xGnb+XVaItFZiKDIpTJymQSjcSnVuTgQbkkj20w
76VWxg37tjQFoVtp9k/mwRVgJGdQz4FWaXaAkvTH0OSnuk4CbO5qcL9UU8aUSShxsGMhdqAOIJPn
VvOp8k2olvK9TufiSt2B9DMzVycp1DHaaBxEXv0SlJtdVUDUSRtX28NgjWslXWW3xbUdkUYB4R4u
0MvMcUwug+QmqWQ6jee90J2aElDie6hklZGNfaY3fXxCnS9Vb8457Z1Is0O5+m7hdwGv/wLthzI3
se9ZCfks1LkWP9VnqB+zeKNgeHyfRWa+z8gzOohh4v9dx/6U22F3eTw58NL/W+aPWyfGx02jq6jK
OZkUxQjGV1PLzP2NDq9eTArBszwMXj8iT2sEQqtRo5NLBequB+gFDCn3aYJA67MN1yAIfYubuO97
vlpEx9r0ikUSOi8bX59m6Hm7ytvOozui0+6eVuRaUUwmq/gs3sY0PtQuePddWiqhdqZJYBGxukhU
x99F4Y9rZwL7x78YjlBtb1CtJynIVXVqeMZwG3Lpvasup7Jy6kWiwEQgQ70px90owklEEJMwy3+L
ETQGgQ9BNo0qIX4MT2hMYrHScSfFjoU3ixVvsWQGSNYhdua1EHhz6k/myQSo03BmMq3NHOuCUMzg
s6ZG6UBSRDYaSWvvAUMjWwyKSsp5ySLcO08H00Wp4Vdq4D/PSBePwVLj4Ml48e3o4jIqCcME5FkK
Y7WDjtevJbDixnAkiqimFPqjAQM6l5zjgHs6Iu4EP5bzAKfYK6GhWkXt8u99jiRBfKo4qZyHeb+q
bPPWtx8TSg54NAn7I0ymcEtR72c46TK3jECsZWQjhlF0I2OmC6b4I5SWAVAxboLF1C+VHOq8YQnu
nGKS15I14/JTXBbsTazr2lKhs2QiMAy/mZ+3dm4wT3XeWyqelBWGrBB0QPP8VaQwng4YjsKSx+gW
QPYrVGJswwaqfEphrdGJkBA8aTYDUMJYvMY/0/dbVZbsRUcBMA0bmvusxaV+OPR34I4XGztlP6L2
3F+vh2gHWBYhp1man3zLEXHVvPRWHVrmIEyWhTpOhFpemA6V9xVTpqJ87m5hZPNxRxi2l02LnP2V
EvVtKe20h7YsYhHq2JH4vahg0Cm+KEEJoVZcrRh8Eayldqi+w05uSVmg6UQNYnMHOT3sUyvYTpk4
hWEAeEywyQ33a87ccFqGEyib/FSYEMhxGnYi29vuseTNB59gFQkqzwZHekk9rE458+UezPRVy5FC
DABkOPo6hcAnnZo9crrwP9u6D+/rEY02NTE2GFELu6dkq4/RAztaotWBYQybggu8qM2Y+KwlRsyB
v86bkD4TsBgOt+yoldL+NWpcJzLlqU6RnQHJ/OPTXC75h+5FRFpuqNBIb5qAjL4ztyzcE/9CJczr
UgJ73dU2DDTVlN+vStrN3JHbshpXpX8VDbp01Vtb3SdGbzla1Hq8d4IMpIOWXkxhSVgddqOPYfqh
gUvu42+jahKLvVU7FAxAP7h2GP6XHDxBGEtuXvsrT0fJRP//6Jh0wMKW67aWr0N38lOp0hlL4Gvn
wMvAApHHKmKyYSY8uFj8KnhC6nCJuu8lCBZEPNFl0JxGMjXC/8zgGky0GnfeFsWqkLcaMB2mYe27
B4Jo4vdOZPUPLPDSl0yDFTAJoI8tysAWnbHSJKA5H43jpABztqnyllsbFoRvoWfLj4hz7WgBTUUE
BgLjrOBIrpgyuO/uXCB/KBwi6zqnh7/MftMw/pRX4soBhZ3UjvHBqBOBn7+DVz/s5jdhTSQVq5Y8
DhhHdAqjoQbFLQBjSrTvwf3Wva6sq7JlOLvCsFbUkfUwszp+pN5W6+ok1WXdqx5/npMpaPSqD3S9
ZM5FVdeGxRKmlZd+8qpMu3a4JF/09xmhLjEy2U6W4gRclxy5Xosqh8I0mZhtMW99rPG7Db0lAuaS
y0E4YvLiXQfAOLTj6H9ViMwvxw5IaMHzLgHP7pjDeERZB4gFkpmW5I5+mUBUtC9C/Qgfs16UEb8l
jqs3YPaSjK0FYnS3/+ucRGjnKimw0nhxhqiSUUvzEtmwlChhuMtfqz79Zjo1kIj8PjPOExHb3Ozg
VFynxk2dCZs3T2akFgZhZW0q2ZwJ0W/ZP5dBC3h6+pWFv68N4USdyQdOV1b8wCdokgaemRZe69WR
J0PzjUvzkgK5xgsIsjGl5p8hFCSv2+JaXY3vOMqjNEWOnHoAUhllXnvo30mEUsduqsh9eQ1lVWUg
WefV1DpAY6STJlO1SIxMCDJqe1TOyy5AHrvIMUPYDPF0ykUxsFYGn8cQJA370h3ZpyRRzEtKNJeG
4YF53JBQi/sLFch3v40SJEyyhffVnPEXypIGPsnRcOgHzLkj7PTa7iXVbYPPckM4KzOQkBHI63JQ
y0W+cCyJxn3hNVHVKIfVEf9s8Kv6OxY/a+5cTAuhCAfvOK3DFzpP1nhaCmHKtRPtP8LYQpR5pLFS
KSEweP+i8Fi2JL6p/MtGw7//vxlf9O5uA2o/mmwuJE81zgIDpyAQc2qIulT0o1kGnYNEnLtfdsGa
nx4sr/ACBxH1t1YrB98iit44GwEglS6qVSBtp18EasSDDSPx8cb87cO3o+3Ys/8efW0SL9e28ig0
ZiELDeqWUHcUQ+gQgj1Xmud1n8+B/eY5j7PvzD9GZUPbFCjljNjyhB6hdT4OcM8iMJ+a52WMgPXd
p23kFy0sulQ69rLOndQw23LQH/83gvF7WyyRiusAxed8tIHKgPPVYxUemsXaXRruiovJf5z4g9gB
sjJYMncbyq3S5XdcDy8RKtKrQDbAW9kXPjOLVO74UPEr6HqOhxG6Z7VRJKqysqbQTaWw1Nn6ckyY
2lHFiQ9d1qWH7jXSHZVsLWKHnyZqIPWdaQngfyzfG/f7Jwek7QZuFDAq0G3VR2kVvfT4suztFkDW
c32V+3WeFU7GSM3iBfZlKcRGkRUbzwri9z/GPvs2/vixXWgyLjeZK+vqu14o6O8o2Lrml5sdAhia
38n0HHKbvxb7XTvTReQxL9D8CyUYQLmfpplBW705tgHxwsAHamiBXFuZS8o+zVmLbGaNdSKm9sPQ
2FRZ3iUsmaN50gcCXQB3LHuCmk80qAExFU1odexuWn3bCQ4gyKNa7XxaMP/jtPrKDyBRxwc7IcMP
QWudlHu62XLh0bf1vW4GTkfGVTQTIqCN+hBMnKBtYQZne6zCeIcxNZWPJ4I+bK7eX1Qn0RbOkFeE
4vj58oGMdrFEXUcZS1tBH9kGLU0twJ6sKHY4lpDLzEZEnKHfp9B+WxklShLD5WzcPxtXZjFqetIs
4TEz5csG2XgCoTVBvSW8V3xsR4QBiMjvxlC0H1FteHl5jc4Up/ilJAs/9J+H+2dUOFt5qjcDy+lq
5zqYTsVb+i3IDrVsMj+BLyCivLHVr2ZNS/BIY8EpSP5bSKS5gPghH5Kx+KH2oJEdDlSqsZxCCGvH
mOuedRyN7GcJydQYKwh6xNY+siG7XAK6ha2QALaxrLB6uBKrZEMwWspvChgkYOWiLd2CT4X9bu3r
RsI9n5MbLH4iQatDf4E5iQMxJz0afmUTrH3iFFHY9Nno+Bc9iqv6V66/QNtIXI3sZXLPwslK4gSv
u7X4z+D5irRr2w99BGPLw3MFN4tG4aGWKypCS+h7hMGDJvMManuhdVYlUNSKU+T9R4UdbgVCxeO4
fale3aH8Jocd8klzIS2uTBDVPPOEs+UW5dd9ArVtM0nf7JRIrdm0jqmGkKQXiboCShlXhkNPGBU7
R3adtrS4TACr7vXKin21dCYdJzcxudewkfL5aTQq457reGkzUVbOQqwctMhx+t13gu6+q0ZuH3Aj
LxZ7v4x9hlnBvRXftwPaZMcFWJtydOW71Oh0tI0oQz66luF5yLKN3zU9QRM6DL6YtAqxOf7qWTcJ
Cl2+sUhpgSCS3zTNIfIOYiLWZET8ubzBPM+j31wSbBV/3z6vUVz4iW7CTYcs6b4ryFjjcglmZ4zV
C79ygWG2HoCsRESZBrYf8xwYnH2ux4n/jc7A7q8RY6XO+UCHqOWqeNquvn+QLv/t7MtYQWLAU6gq
Kz1lscH/S0Y5D9UoEQCu8r34qi4Ah69PpTyN4Q6YdpeVIStwOKlcRL2hryqUvUG5Iv/XsgkOnzw+
WXFu84C8fDQBVEuP4c87Du8qzXrKUfZCn/mqXJkHZld2lsz+C29SCOO1Xvc4J0nQWn7uFcfD0xa4
6h8BY0XWcl5PFB+wvhJKzgJr7H2dUYaiRfFCM/kEDJf2XPcTxTep7UlryzbX5FRbJBZJEtn+NE0w
7nb5ADti4bsnO6zb8W/WYKeomGTfr6uki8RUDEl2ztTQBm1j89JxENdeO+wLJDqT+wMWrBrHIXTn
mmTJhv+jroBNmiMu2zLIVB874bgFm7q4Em7xWBXF5WXUEl1DuR5KZOmh0V4N+8F7V2yPtPhk38n+
OhK79G9mxHQuIE/V9wmvFiH5M7F8dYMR/obPl3K4roZseSVoD1G3ENCxNsA65Kt+XYpP66jJ1Plp
WJAnbw3/+z1IHKtngaD59i0CeBr1RaJB/wkOyuCxDf1IwoNP1ujSzr5lZ59w6X9CdWv8QMZzHQ0o
LG2onYq4tYqQ3loEHER9ZuW8wvZjd9qVqUFR8fdVQUDqI6BAdXig7/R6/bRSN6KtIqB6dKPKmY/+
P1IQrnRXLDFOvdgaOxWeZbeCOWuxLje/x7vBV+RMnMxurZ+Nzy8tFPSp8SmgFaIcvdHG9P6PXHub
cEauVThNIh/+rIOwioYBypwq2O2ii+PHLwtLmhucINE04ta3g7zoRl4s5b3Rz2OIyJbQxPrBmvUc
ooHi476lc7q0h5Z4VajY+XUDD1sbRpew/7F1ynyco7UmMuaF0GF/VThpmEu+DlJRHbIbM8lf7aAI
LNku+CVglhv7JKGM4g9oCV1WHD2JPWSeQayyp0iOyrhNvLrfIP8WkknsLKbavKjBaT49CKdm+5cp
X9/ioLugmWZhDNOSbuGtMO/lX8naZ5U1qIg+CKVaHPpCZ/u9Vq5uRU73fusOTo4jl9ayBgtJ/Qr5
Ed81IiAdc1ZBKS7jBP9Mc98MdWxSYrD5XfwfteMuwwy9KfUFRkS+TCBW4UBMdt/ALhatwi59VU3V
tLhkkMaYTyHwnbDvL+iP3LHWf/DQLTH6Ph3gtrwhH8zal624bKowIQC+yo/peI5AwaBWdf2H2x84
Vb9z8Udd4ceNtIPTyrI8V/bvFQ/GPg+uFzliXdBsWJP8whr03YRal1rBLhYJDpFYX2ge+QYHEPZ2
FMqg2695z3SvxLQSt8+4h2adgvYYdBOFLatonUM7lYVJczBQE+bJ4NorCwRLS5Ut/wB4Q/ZDpO8+
F7YuqqP7MsDJPbmDElJqxFQ+HmjB6rEgy6JNfTfqcQTCC5elOHdtpaIDIG8RKacqffRtV0D9iBXI
c7DrQDJNV/ueQijqb12/imKSdC2mGyja3WbmmfM7ONI1pW914ZCg0CnqTuNtNiS8GheYN7V/lq5h
l81VOcfuNrIJcBVyDftL059nJ1RxxQNU0JgygAuMvTv5N2b0M+Ch+CYTm8vT2wLLVBEr0QH+eYgS
YB7H8c2E8FfBl+oh77PfCYJdEEBqPoLcqX1yjcSt5lN97Qtc+wyF5uxmWV1EQ3N3GNuLbn+R4OKh
mml5vX/5/MmO9fEBKp/luJJ2FRyCvpiDEAW6CdH+7RXgdbHXdkGlDUag0Y9ItNIcz+CiE8Qgmi+f
ApS3C+x8GgoZ3zFifPeNG4kQ4oY8jqDpjM+68MHhAcwQfxJarrQvrrbKbPIykytIrm1poqHGXt/b
KeRI85+RhG65uBPX1+F+55d//e7yqBdUjVRumvXHLlSKmrj7BlPk/FkmuEQ6DTpBH/DLzUGUVS5I
KMoqHXeLWDsOWDHLPxuptnQRxgKuvqlkB4yecJhtUSaNay8xBT0eGvzYAu0HXQvuGDRPi28CNSYP
QqDt0zk/j1WswlQrLRtg5VjgTVj9itjgj7wtcObw9dWGEAxk44Y9jUGuhBbE/w4aP2iI9Hto3eoE
xVEH3kRE+b2UnNdJpBA6tnnkmSHVN/BN8nlef86cmy75wVCai3dPFjbArEFfvHyPesu6ifiM+D3s
tG8U+F5q/dlzmixdiwrhec4V4ND4WlLnXMSRF/0672Z/BKQfhpjdXSz6IYPvX2dFwe0rzEUj+s4V
VqlMEFxtySLsgX83ICBHEmeyHbklLBWesCuUci5xMwDdgRbVErWccHExQbpfg0CyAa2YUov62v+2
I9dUMTdz+2XGysobIkvNptcWQ6R/9vxINTQM93Av51sI0UEs7flqzuv5zVu1wtURM4HNKRgjYKh8
1xXkHHUJqT1NJ265DgKhNlFI8FBfLsDBNoIcTUAYpVn/tpcm8LvfqE9+kf3Tb7tWrJ4OYb3jUm4v
QFDwaBIWO1BJWZXLL4ZLrm0qwpIi1s70Mzpa0O+hFPLfRPpz98FG9TdZYJaLzn9/br5k2ELDJrxE
/XSuj4uEaibvEECzJJXKnsezHbosKRGmNxlNlhPQRGXfba7ogOQKbR1kCpfYtG96UgSYnyZYPgcE
qzJ3QcVpt4dwUsGlVCA9PSpvJiGmyBbwrAgZ6/i3b78RXazUWRrml5J5048eulb/lIYM5tLSVtri
4i6WfniSzvWrIOIrl7qO/FopKzkFIjDx9a9t8pnqhfHb1iPcwGPfWdSV8WLFzDmqZ8kiDUWK2h0/
aKYxexOYq3xHY2jeDimTD7DW2f6SuLCFezzl5WVucYyCeUzKDoEtK95s6N7R6noy2LHYEvkvUvFf
1zXXy0OdTWQN/dK80MukY0+NlEQ4vmXuo6j52UFlvVSqBwAEihNnnfHKtBSX1bxcmDfyNdKoYlLw
Ou7VIoGuXytskmo/D8S+66K5V3WjsFfrJ0cagyQDd7hqAoCOeQgGb19G9uWhhvt6cuMXaOee66Kz
LtBSfL9lkvgJVv4DBkw/pqXi5maKbcvJyWLtSI77FrBdB0Y3Ek2+Q5IXGAHLvlQEbKx63GXWb8Nd
sb+LDrXq1bawWxUU4Ioyuy/tU+VvgMxuPuUQbLZGzC12DnMvGmMVB8KUMhvYRphYqOcMrSs3F+7a
iTkPK+GUP9mkrR7CVNiuX13oRdTBY2L6MCkxr/3KiUiUzFqU+02G3pdH1fdrvgTn4HmVnq9Is541
kqlCeWPyKSdQ9sKgdsrcGu5EvjBwErKsCADKJfFM9KuVjP2ECKwkW3nVN84dbUjXl3MGay+Yp3QD
3Ql9CTO3FCnQJ2KDAq1zEnxaO459+Dl3Hhe2zHvdgEXdsiunWdAI5+U2T89dBekFxyC2tAbWjK2o
pxIR/wldNm8KE87OAM1axdZYfXgIay4MJstW1U4qj239J6TYVbzdnb6m2VfA32Oi4hmueEBP5lA/
cNh8fx4af7W+OO5Fd7Lxew3K6FXd2djFvrTBRYuzzLmv9jCMORYkHbo9j9ylk+OBpzsPBDqsBNjg
dPd8M9agPa66KaaMM91FE+IFp2oBdaH77eF/1FnLW8zfylZ8OGEbFtKR4Ihnjqx73j0vFt2Wbgy2
M8CQROP8bXn1d6zC7z5P/z54ko527u7BUf+6zBKmZNZ0Yn5hDrO9CjzSyKGPo+FI5Tu7Q3sdmKTS
w6LmaI0g6HDTpUSc0xHswM2O1RQ1CvM6iTtp0kEFWUsalD/hAdm+D8XRymsk0pF7eo9AqSlYcCBP
2mOZKV2GEHx8qfE3B6IK3qmbb7fynNwQtfPT7bwtnq6iDDW1A+YyRZ2I6jkzzbE9wcuawm6JrHKX
aIZD8ENRFAr9VIlwqf/KisB67to3die9jsdRk17vUR9GLYRDBIPlIZTriIdLpaArDFXEQ5tY+jfn
fk/its1l11f3CQ2SIW6O/qMt+ampOiOVMMtSjdvhcBfWzBL4nF7YcuTCaBr0tJBcKdylP/Z1m9t5
kWZpE8JSWAVVT2y6nYt9UPAU8g+qt/yhBOy6bnfslGQrofzOeFa8Mr2VhCcjtwBKOfmWdOGOFEep
D3I0UgTuFqx6Cyiaj0syBNUCjl2ipGKKldE3hcWTHIWVo5n/VQg37pCiVHQkkQPfW0HFtshM06sw
yNYhWt1etSaIALuuMONmInPIUBT2FyXmkIPnKokPheAmu2b89GKY/CCGvQAPdHH92KB/Pop7FlA5
OjqbAUdGj2HpltnQMINyieHETJO4TCgMxbrRwHkp6UNNBe8u6qUjYXogZNtA3RMf58S1pu5exof0
ttgwJOuzCrjQh3yotMT8XVOEgrnovNNdg8mZnPizw4FwHA7eUJnf8q5IWk/0uR2nsdcF4UCbk5vN
gcvf5I4iwr+9IEnKL1qFqb29+ac6DH410aGQ1JL995I5KvTBoYDqIcMQ5bT93LbgXX0S26KEtlCa
LPP3xliCpc3WX/2kWIpP19Tpj4IF78rXovqhk5gabEycxOB7+y9pu7p43k9vnGXpuoST+tN1So6C
U5GhWMxsczU1O35JAO6XePOaloxS7x3Z7KIwgFqtRKXiJlH9yhl2yeGUMA7sfnrHZBlGE1SZjpeW
8eybRxmr73ghqbAYwJkngTfj0iyCgBWYN9f3Z2XRG1o5eCecFPPFTvMu58Li2ykagydpArTNa3k6
JX8CEIVr99g7pWeHaB0ABt8Jre7lTjTXj3ocDMQ7HozjIxXSjJd2Ag0+3ZnUfmGiSDLCj8HplaMJ
+7Hw0GnSZ5KC1fhyDtEWFFSYs8IV4oZWqtOplXAa2rkVaqg7TyeUJJ6GanPQoNqUYqPGvbNN8PSK
oO5CSqnqWITvvCyEnp4afqmy6610K0YfQrHMj8Ps7XBKTC25T2OZtgrc9wVi8zS9oUGUvOlA/Tya
jumtAUnEW7QRtcjnNHToRrHfNbAloLQBw6EXRrJvphbg08LZKmdjc8rvcvPoBpXSJ7Dev2tQdlSZ
DxoErIAw/UibXawgpzmoX6lAuhb27GKYk8Kgf8CRYlJN6HV0dHel2kloUxdw5PECLCXER6oyposr
QuKlg5dQFjwAUvwcJonwIEUchWvnDEg0c9QCGq4DOxSBCZfiGsTFbIyXGGTJBS6JRr8cGjzUvgDz
kn3rKxhnZ46c6HCYtbSrhEKYOlEtXRV3LNfFUQg9f3+tEE9F8Q/sSGn/0y8g+cDBLceyzfPx2esB
znx8NAo+H/xz+I19pFy5FwjYFzjZdpZnV1nsTWSHswixQUaZ9lB+3fMXcPa06PqDAAAzLFVhkA16
RSlBnF6TyCJ0VSb4Q3NIb78orprnXM6JhIeeBJbW9ofyybvviZPM3WBQfKp0kAbd/bbvmty7odPS
rN1i7Y1yXFl5qrRdRpAzOe9dBi2ViCAbI08XYOI7ZOpwg7Gml+52cucgfFlHiIvCLrikVnpwp/uK
g4a25GIH9w3CBEL4nqtwK7X+27DaRFmNDcoY1B4OmNwHreMrMauGh+vORG/Xf8ITDmz+j4GGP0UI
0neqWVPFpixZn/2s+kX0lWvhNdpkgNF38yTLztVYOmmVy1SAayi7yuRS24sztqmmzJBl+kj6GBjT
FWWFdHeFAx2bCcvauwmeh2B/vmoonI/kgzMSebkmgULaVe8PlxhMpJWbFn4PLi2jw5eoz3MSX9EB
BAu+VNQGj4zCeSmMTgGozqSWwqFc+1jKw7x9D5flX0NHwI2zHsqoqUwzffPj49UXnShpgz2tX+8k
rK1FtVQLAWcFpvvwYQ95Hg+KvlCCsFMSzWNBRzIWP6EZ4aj730fUSnIV2cPkxlxVMZMhJv8gpWkw
oGYmBYf5Tze4dKc6GYwTIyl3xHP7rm+4i/h0zf+Gv6nWKAcJdsv7AvL/qsh+rONy8vi5rYRkwPQW
y3e4f1a2ONFVF58NdfgNC7CnkEqHGOHj2GJYYA8SC3W66aUB/HiQq+B61dExlInXzps3dS1B/E1x
Wny2kNtmEicQpLe0E+yicOGnymdtc104GEzwFcH2hqWg3nMwxXCYj2iIghzm15DPg2ZbOwEgyjLo
Px7qjKGAphFUraUsIsJmNFrHjpRFRQ18D/0fnaDjD1TDIrtUx43XAY3BijyGtQ4VD+HYSqFXT1Jr
whWBP3ppDvgd3WaH4xb2P8I3zmBUQKxyzApQPEMCSSSRcYmcIbkm6Z9vT+yrZUdSWtHi0BlQUj2/
yJAGOB/BpEEaonWGhsziJzTT0UQq25ZhMBrXI4meBAYrtLfki8ym0spzkOqSMgyQL0WkcZ+Uw6N5
8JKvUyVIAqCqQeBwKB01GzfbdHpXdKhf+wXvnyJkPtALLXLFo7zb9tfwf7kzhRDEWq8K/QLlfMZb
8K3E11LuG3PXk2IOVXemVVjE5H/9X8VjcroGZL6ybRS+D49BNquJkh9GjyYTa/kku8uBO4O61zye
x5+D8bg8bUCqIGHmA2RT3cHcBNWDqgfiKhJzw6Dmdv6ZCgt2DZ9vXCWRY4At/sVRYQGAjVcU0LJL
BRR3avGDIH8EijWnRua0TuIRPrBWsiVeWgeiiF43pOlllys05QMssyK5B7JdW+0g6Im8pRPo75Ni
FWMcarDnW8VB62zYlTRmzRDqyaCNRjuDPRxNqM4Uuvz4YipTPNqZddKa0jTaHFj1P0OxUE5+rGEw
h0V1OKmQDhQ++i690TpNrIklQqRPKm7u1h0DLJPccQW7mggiCrL6ALzFmAfWyTKWAKTb0CssrbVd
Wt9owzDQL6HWle/31jhdqTN3/L3kQHYbmgIpgCqb92Ir7Myae627toZ4/+uKnDX42tyeIyjfrkz6
aIOhzXbZoMzZdxWoCaM0pM6A2y0JOvCHWD6eO4GBGeAuEtDd7ubD/roIRNutxb9ZGzxABJz//sli
fJZ+U7+/Ra+hhpvLhC78Yy+kionWnWeBxfELmPHbzVwiPntxuOGY1s+xMZvX2inL+pUxu0nUb2P7
LVMMF5uzTqqfvC7Nvvpv6N7YnxQw18dOEgqb23EbsRK/3h7yTul5G1+lgtUP3Q4Wf7JfhN0H+9kl
4yTYuQ/i+O79Vp6lVOoGRry7RObYtiI2iy6EQ6dy+NKCmGEKWcquM4e5hSvctdCQRzqosacUdUYb
JVR5FaWExBRNiXY/IxxQl+EjyeadEif3+E2AJW5Yw9mWiuCy/yPT2SvdVSAV3mkU4F5Ux94ljNqu
7VoPBZ3ktIHsz9GnV7mxkfQtp2cNH8iYj//11ypsAi/NEBxzGCkdtgP6COQZXrc22ZFc0RedanaX
2mQ0xvKxPCzUy/28TfnkWyTcj3TKQA9pDOeaCZLXazGBZfZnbvDx2JLfRKjGu8ZUIHVLsdV73/ua
PhyP9EwU/A3yzIST+4jbPD9RBhcW3yi/7RLk2o/femacLwhdTCJ6jtjHlPbtWqqRmcbzH45fFvTC
bVXy7/PvIw3YhhcuJujDVZQPNAFQWUXfeZBaCdHfbMmrUGlxnyEaimHVljEox0U10Ixv/99MLvlZ
eH6IfSg9ocs/gI0qY1VP84szvQ3boxKOtTadpdjXm+SA9/buigw07fMdt5uIVk8imZIxLjEig91l
/zGmqVcoPRvpSpqG7j4vMk0XjryFx2rl4aaIHkq9yetBPDV0uMow9lKVEYtZoXbydV2DalRuO0fV
X3nauQ2zaw6ZredDpsnzEBREvT612h6ATtHjJeW4izFcxkqPYs5Mmtc3SttBib3R9kXLDA4LL6xD
J3ectP7BnMf/xf4fB30dbjAVVpTFTXO1qK+gcSBCrZJ2qULDkBqZBtML0rauWep35pD6GpIHj2vh
Aar/eggp3cQYV85iyefpUsQ37JL1kms4/Cw+Qv9o7ip8DA6AwAKBW9e7ODWECwLlcXZoWiSWTfQ6
nqR2njCzjWMDQk7EBMHg+19B0mAjwc54+7gcFlcWl2wJVcEk6dDFvj7fk1MV86l+L4PFqngYrp1W
fClULyeWAAquDKZ3BQ+Y3CimOm6l3E+TGxSUo3rbXnEyJJsWbHfoRhmQXsg0GwSIc4hNX0c9Co0u
vupSD+WulkPAYYciqykoD7EgLC90VgY9B0fySqUCS1UE0oWg95/Tf7QuCEEpaOvG37H+5eZ2v8dx
Js5+pv/lMLyXRe+kkPld4XEZ0HRDYg2TAqFE5itLh0qUWbqKPbFEB17NCFBhvD4wnsMmDW1IQeXJ
5VYVtW7OtDMNHgiyhof5OAI9rDAPLXvBpSTIXgWLO4oRmHifb4hYXR7XgwvYmX/jlEAkUb7YsBZx
bprmrZ8QbNq67EOGsVPxFc/Oz63ifLannQ5DV1jyHhi7pZAq+2lveGYqzRgQ835oTxjqr8JcKZz0
1FYTuulYf6GuFOKEnC/v6INFv3n1+pL0+S2GJzjaxNqvfzvUX9nX52B/8jZ5qHNT7DMOl2a0bYzC
Kkgr+th1pZ4b2n5xAnWR4G+tgav4jvVbbgCoD0jPoxeDZQS628/jo86unUwv/i+ile6n/4SFLMZS
lHGnjp2NHYZsuihj0RK0eIQNyvMow9e5PLKmXAxiI6XFduKkHFHk2Ylk17BgmeIO2f0rW/ef96ds
aIDLEOEDHNrkb4J6LnYwdo65w/DC3wMVLn8CCgJg5y6MG/e/GtqKwQ/3VQys7zynDh+O9pVwCypD
YA+5Wol6nJ6smjbd7OBec0mctsWs2UtyvBhYKw375BA93ud7Vk3x9jKjaCotJ8PaG9bzXvY9hjcV
limcXOlbHPErdIrD4ZRWCGVh+w9305AskPF2szRWe61JkWNXn0KHAmnz5+2cSXfQ+UizLiMPicpS
L2UUR7YSbtKTsJpefgQ5JpX5e2AmMp/LGdyqfiddLZSSFRd3Mx3t1b6hAIYJyxUk16UckASOH0JN
BlL4OQX/+5t4ucHPfWr0fmNWmbW/v/j+BOs8ZY+KS6zCwix8j6z1gvDAk+3KeCBhlQ7ou5HepLsr
DQAkzxw1OAyN4PTzEUMQuhjRn6kdP5yzMMzLPJnD8vq4TALB4JySHmVN6kW6f4vBw6etz3omFPAQ
uW3VT/NsiDBmS+k3hX8yMvxqnLAVMfiVts9c169/p+SpmupWW8etOtaIq6WfxqLgcnWS1H+8kE+Z
wfOuUC7z4bjy4m8i/gsWoeqnhsmc+r1xirbYIZ/iOeukEuHRV7vHLlqONkVx2a8Fgl89cuC+7oEP
VICxrFvtR6RpoJbhxbyMumDjJukDADRQDP66u5QiaBtEv3sldOfu8CaHNFAS88uuBeuO1WVEyxT1
80/t0hd0swiFJNLq6VuN8ffDD7nCgWjZSrenubZDQXkqfdxaA3iOOx8zmSOC9S+c6xq1XdkctZ2Z
7zeMOTOTWG1AdU2DWxW76ZaFSY1Pl63ExRwuXxhy72kWq5w+c2zkob+UY9edi6rIhrp/dK1f+yYL
xDAe8Z+N2A3Jd5JTFhdxwxk0iKtaayKVa51nojN25+dNjJH7H3ZCAvRPIaOBCyT4Ge9Opg8y6ct6
7mTN8yPmrPg33HatUa5u2C/i8ife/RoFPIAq6NUEUxcx6THzSAVywUSd0FszWH3bB2nQeEdFZtHR
LbZJnXWQwrb3NyJgxSNfkmxJHwtygzeMVN14RXkIzVLZc5TNH+LcbX6xKCMNjqEet1AF9pNlzhWX
cii2o3KQWr8rsrcvHMzWpLHApxkh/Jm6rcDgh29Dv2jdbEtNBUnvxVFrZlVB6GcH6jWsxk3cJWkq
w8GrvjpRwzLhXboD+1ILGlM/LQ6xb/P6jFHsVdZ8Z/sgKlLGQMNR+5Shm5dU/QQmV06aCj2MpNDp
JE8U1T1v909dJ6XXBgW2T4qnIk08o285ZxKS9D6ASHpx76cTA1FBEKhQuwoero0ENZWdH73yMvgF
R6/BWg/XuI462JWT2cC2ZSaS09gLCixkYwXZM1KCl2EpLhnc2/ySaHrMBWCJqSu0Np9OHa0knsOE
y26N3zwp2ccfl3zlnSP1ql7VCqYQGtgIDo3YIg6M4zpjqkhQsCaynYEtyIETEd7y/5+WptS0BRJy
PqWE0Rm5rrBo2sc9nKnjNHRee/EszYn8XVrawEe4wtWlO3ny/BkHIBrHpCtSUyxYB4OD/hNXFYu8
z6+dLgt8oyt13nSxxjIMBrzIfUTNoQ8E26+VOpJSLoljOvGh5CvsuAw/x5UemXfjz5vgIUqdhh8K
oukQ8bhIixwpJBrC5Kdy/F5ys/vskDJ20gPcaClyY2xLgT7v014f8riICcmdkIO/kpTSXGTdBvsK
b8b8rIIPf28fKzNxy6e3+D2dNqo9g6I27ZDnCV/Ly0VhVB7nEG007XaGhkr/aqK2RFilnTfELJFl
jjsHqZ4bSZj6Xsj8yS7OOU0TRiuI/MAYOMwBkhN1KknPy96vkQ0ON6F8/Pq0OXddmjWTVuPyP4LR
SsF46E90Fw0d9xeu1wH38Dkcn+xkZC9whPZ01qo2wJ182+Pv4lTC3hwEBIv1zgq6wDkwgton4+nV
+WVwYA+rBXAixzk/ZTrtgcpSADCNxa5xIXnXg3oIVRS3qsoMu7/9jMGC4/e6esdFPR4ec6oA3cFq
i0AQ/6eZbVTs5WmveFiBGz9IAidJQ0PNFrHZKu55+BCbHPXmT/KEMsqN96h0M9LG+59A1pZpfg8C
SADvEuTf4BOD38FQHKX3vc2/feyCzHm0vN53ho0Pi5E/YWPbZvv14aT3AVSHbxtSMjAFpQ7LF365
DkRKXRFtoXXXiJii1298cS5pAOn/SpJokeLZlOWPA1sh8W483Ts6EEOlqCaATpxpIN+ckjZ9f4Yn
tohJh0gYuKp1+5DIzue+3btXSCP+PUl11Rw/Npd0ImHmV6xNI5zXnCzrgIXwJC6MMrKUkJRBr9CB
uW5E2NbLtxlgLTjt/FJfYCljL3uhyDYWTAsDbA4gh5Yt4vYUMTuHpJy5mhzNESZTuPvUyWlpv5vQ
FtNM9aa6VA99r7Vh9xu69SycLbPtzJFLjjT0Yac1NU0+A1H/OSn9+6AP5yPw8oDxK3EdWDeBXJYP
entCkOxhn+aMfRVecz0PbPnm4p/5DOVcFETsVddECCGcOumTwvPN62XEcblLsoJiRfrBsYhdlHYv
UXlgoSrel/9a/UZKrXEtL1zvko9+S6h/ElrMsl+gGg3mz2A0VOalvVuJp75aoH1uOF1mahxTDVId
Xpjs1WnuKJ8Py0kMbS1rXRjdan4+s9g3hPBMAHn3T3XwZeIqjGMcC+Mf4LFaCfx0vhCfk/cpRU5o
DCxuggacxak42mA+8XEh23N/H/TGvJi3KGwVTW44/g4pe7wK2rDtzOZSDAHktTxdS1wYS4awBBKz
CHOOVyzDL9aPOYGbVJsfJzRhspKrxtDQ/20P85J8QqJfgsP4RNxCCPtybbgcyZuIHTZCPg4cbKIE
v9YfJRTxF8t0YG96SkaAaDq0xuMGsi0TyWNsjqEW9fNvKUCOKg6oI70b8uZbceRPzxmVatTFveb9
sTn4SuQ+2YJi3D51B9Fb9/LFGAFzh+m1+rfRPFH7JJ3ELp7+gf/qmnGzCsCmO8r2cMDaFLb647f0
h9dNLjoF9/jEK4P29xfu6+Ylx8VshAkPn3pbtokhFA6wlIQe3vK3MXm5JAR9uDzqsh0X5R12DNz2
TwB8a1rmZOagUPUzKcPUsOXEstS0hoRjBJKTUp99JpPDihcM+jDUpfmVSuZAbJ9BYKIHLvWaSiVO
ao4QPp2aulPSAAtyIsmEplLZaOEefrqAF8YgqDdWdXbxPrcaFF1xUZNZBwWFUOQLwqGHFKTZ+HLC
eF/shgk268zEFCkrLA4cCZIEGv/vkEVPReTWwV2V0sub0ufc+JzpjnW+bDT7eLYqAZJ8hUGJgKcc
DqdF+kR1Kvma27yji33vzEQXvOcLbpdZ4Q4ERRpJ0RZUPusuKJWRe3pU4wuwTPh7nH7BQHy7oIuf
W6TWuibkr03TCuYxkycTEhti0tJGGbshcpLdYE19Exh4zOQbhx9AVoq/6djalklA48NzwbLjH4mr
wXENcR/pK0aMnM/qm1bQDd4uSWgAFfE3Dey7bJxmOhfMLJ6UtdP43eb6w4ihl2vebehZOeO8hi4K
7+rQQ7Wi/cKeHztxstRMr7PNWFIjVid0yjfjEGzdVhQ1StcmihgmO5kuOta+7svf/mDaScqjzoaD
FVeJBZuLZ4zRCcvABvelwidDwHVN15/TmmS+Z3vMWF8vqs6+ihm5R8vSGLyND4/ERbAxhZawyNjC
b7ejKZwZ2nTKV8NEcoeWfsSIoL2dROSj3NAbBuYWGdS03A2r2LlAPtBCmpQzfrEORFOhiU07pCgb
Ewkygx6EQHEk6FpvQdkqBLdkX4YIdlXduwIsWCHJjjCJYZnxruOGAWxBOZRN+prpsFAgtM/bMj2U
2EmWHC8c9EU/bgn5wtv28zdQ4BAReFZKW/OIU4mY5CPcW7AQ56oAGLLijTKX8L5HkfhmMABEQc7E
9YqucYAfesHoGElEHlCnmdpm5T7ed353m3tmVNwRJG8lDwIXHI3Jy34PRUkfs6R/XdNW8y2vFSbH
YLOS9bIyHLnul24tJuHYa246DosL5Er20rZ3VZiQCpBIYYRBiBQA0FmW0SMMi5ka97D9Jv8UdtDR
4Et/XkcNpxwBBg3LdNHEiRGTo5jhB37olz66at4WM748bW/j376slK/V2QxlmvFuwM44wxdWnlex
icHDcu4zbuerWiVncNh5H4duA+8/PWwIh0XcEUkK/QwRVd7lzfr1wq6Arv5PSqtYeQsTMmcrcs0+
ea5AMHGGybTReHKM3VPrYM8FbshUHtJ/youYCC2ebpTNpTrPe07gOsvvytOje2dps175ZeozCCJN
xvJrJvYt1Kys6ArSoJwjQWFFKXjJ8O12BaWpTVhRRQNY36UhaeJsfyTtP1OMCedLApIgZ9O3QW6G
MbnADkKxUM81pGJt7usv/WIwJ3PiAMvs0ZBpf7TCVHQh1MP5lNVd3cQQKXQl2gEB0lTY0b38O1Ay
Fxh4mS65BamnBQ9VsGZUN9SwR4PyorPOnXwtJiZnC76aaBPtMZwhtm035ByzcLNAV91wUH5OPthn
DH7fW5xkGdmTp8xPRr8Meii+6rVoTKkYMqWvpoZw9PY2hs1l13xeYfzEEMeI6xHrkJyC9gixXyby
sgm/+aSSW5fScjB1qi3ORiwf4rjOhjb2W3v8UR+K5cWE+81GFzVK4T94ggOFprPiGjHDUj1cI7S1
fp90lXpk4stsQPGmSLWXabyvNheT0NPZmS4rVGMyxqAMwXVqhIRS6bYbAqfsDl0dL/aFP1MmqG4t
kNZuGOLuBE18GojRJwglJkV7ZrJVc8tKc+T4NtciGeFgrmsCO9UJPkDLKGjlBC7q+7EKflZWF7rr
+pBDy6Q7s8saV0g2DnGhwQShAbjHkLea3l0v4q+vUblT6+DAQnptdLFgECTLTMUE1PMhoWwzBxwS
Vpxun1vAvIahW9+Jr4BOdVJum86peMyVTWPieEJHq/GG0fOSMEL/cVdLlAE1m/uKqNQ4On+dB6Gn
o873hn8G7/vjEtkd6pcVRW3Igp/Ir8TUHT0MmqsKFg0oRrcgLT5ghKGCGTMe5vvCcFgGDcd5un7M
ZeIrolYD40MIJ2V4YSVPX57Rtt+lXJwQeo0wYzANis3mdt+5Abu+Vks1L5Y5yw2hwBDjHoIvuXKp
76W2VMx/rLAQPI9FWAV2afU8IOw/sJaeQkp/0Va/0CuG0GMD5TgfnlKnP1gok3K8UaaH4MXz7eav
gv36mfOP1Fgo2JkxEBoPqPIqE8qP7is2W0+zJOY7gxuGibCxGcYQQJ5e/L2jR5JTxoz52HLj7aVD
CMNRNW3goHdOJ6vHJZsy/DXIsIcwcsxPnZ1mu2S1FffICtm3qdHZiMYDXraURBbgu3IsmPEGdFLz
VwanQmZfre+2A0jKMax+xlt6uDgp4zSqmU0Tsz6ZfV2Qol5Kr5nKD5Q26qRXhLCKXOhyFhXQhYQo
r9Zay8iSoZP8rV7gdb1tMxLitNiDYYnyM4ayfcedg8BwCAkvFe7moKVyk16uCGvfduXeRrA/22zp
vDslO9ySWGqI0TJw4jrw9YC0KglIKSHO8bP28918a8G0YFUGVtO6FG4CLpnMkHgg8hleDvCZRWCS
Zr4cJEFtJHJlYFYhfPMCpkbbF+g0On1ovtl58tV5eyh+dpetaxFpvMt3EPxgw6w4H3IZ2RpK9eT0
+YPne8DZS/Z7AAGcKZ/ubwQuqlXrJs6AsoHrhq4iAWh/oy1jrwtUMnz/9rq8d3P63nPdSe1BXoay
wRX3wK4i6SfuRVp7o7mrcCsjVdKPLDePlvSmPeLCQejQrrFYQxfqD/0LeXaPL8rOEq/Kb4keOTS8
1dIIx6DGV5U2ZS/2MTXWuf3Ikmruobx9HznbTRzG4osCaYlFFw7HZsxPgT4oSjV4Ufi99Q65XpQb
rcTgrCwxPDCVnUdgzooUwaIZVN0gmQjp8h4RZzBQc6xaAfQs/Sv/3JNz/B+tcjfu6QnM+EnsxkE7
fx4j9KRotNJzk/XK58XAQ02+fz9T5i376hARk34gYgTVITkgYrrBZmjLdFoq00NoKUcgti0VXoyq
jcW8SCSjM2BZszpkwpwfMYzLg1srl+dYoO0RLckDETNknfTw4TkwcZdjlXfw6j2P6LeFVRJAEdhg
ggTglPOK+r9/svcOeMqZ3MTSB1cCMKoDgonKiyf7hEDPHDmgFpWjTOjRj+CLF/jwXz+jZxZyTx86
nflpSEV6QBShvVs3y/k022bcBhb365kmq9JoSa7JNO4izey+g5V7VVGgTU09BZWZuedjBIfcWmcO
8kGB6WLSe2Cj4HXT+SDIrNaFQJozKNnLBIF6CcesDbgM9k6zgrLFRfOSDpFXvPzKi+ekpoBIamg/
jciRKY3a7fZ6u/QHYIu4mOo0dA/1vxmGxDp3AUT+d7y/T8DBS0PSKouOLyIRanmq7E3x2bD9KR+v
yPj9HbFnwOyZYGd6CoNzo6OyUqu+EQ+jOQdx1FOTF9hZMhMq+RQ3X+rlx+sbnJdEce/zv7OaOPyl
0bggCGi6X5K1F22iAuhSFZKq8pj8oWY/GUkgkJphvyBMu3YPlQLnS3tef30mNF9WEDbK7QmkjMmN
wvHdZXwKqPrqHNf7/9nkg4MPww00fGLW/NZnVREy0XiPTzAOpMdXNgyetcu3Q/JGN6WsItyTxFN7
jfXZOHN16OvAT1zDDk+HXLDPvgNCivDmK8f13LNybPlmE6v64blTjwAe3Z2r6CBAvKRhfTh4P7QQ
C3ZH3ApJoHfoDl4DcqOB3eBIYk8/9zhrbNM7kXtWph4u+1KLRaIHiFmyFzA5T0mTq1xiTToZWCVA
kZDh59uXfUEEKgWTDIvewMatAvPdTPga0nWWQdfRvQ4CLmPMW5jEu1IWY9drR0YYQjjQhYHnNBnq
9NLkT4+1+VDE7kfqsnrq/CqKtTefprl8JR6dKxzR8ngAYOp1acvyaaCcXiZIncTlIr3bXwFlqPzW
ELG5XPAeFhDHe8TdaoA4keBHBc3RZtmgTjUE6I2sAhX7aB1GH45aTS/2NsjWhemfk8t6zQ5w+vXp
s2IPsdd5pXxfMSYvOsQda2svuHUy7dJc47DRv9KLdtIW0REIAIxPae4+3vNO6S5tVAZpOb3vMChS
cHnALV52HlSl63YPFKVAVhH6S4GL2fAb3bN7EboaYsDhPRrRrgGNcZ6meUkEgSAK2EGh+MDspVu4
l19bULGeleVAIG3hqc0BXWRP6iqwQ2dwMeySDKWpd6xpYnSPd0wdXJHrHGART6dGkS9iX6Uruukj
WusYMwU/nXFeO6Of9AprbMwjylSxdnK0EZux4+DIS47xcDL1yoX2ZkXJ12Cg6KUUz8jHT6SpHdT4
6Z5feKtpK/ywIj4t9ofOUEAkgiQ7U/xpZbOrX4byZjEeDRJJ/R9GYnUBjHrIzvWJOLdzHPcp/yGH
owll1zjFQvyzpYCO7CnbZczxUxu9nq56CuYzjoOA+lcT78uCMvffzoKN/GLs697DVde8e9pmRQvT
WAv3U8Qg+DMFK0HcU/P4CbMmUB8yhavto0L+uC9CzFXfHS8Rp1sXkFzr2q5SI2cMsk1g8RVbdJDy
CheGAM4yJP/qH5kJgQxh6feNMeUrJxLOhlx8Ph6JsgGwQVH45mbDKs4BFUHpSdBds/++R8XDQkTw
SIdiHXWysRrRx1R1tUzNPLQH/U29wma/G2ZSZqCtDn+53nXJswd8ZhtjbN912MDyHEgLka6Wj0Os
uI59P99NCzb0YKqH/TjibWoNFBiBK7qHYBRsJ/gbp9owNwwmAZY201oa1FM+OsP2kJGEQkDZM0bk
s2pWtWzMfCbhW0JFln0zX2B7gM04KMRJkdtdpPRkbjuiijynKkccKwQvVrr3u/tqGjPI/DzuNUdk
0AN2eVUqa8l43JQim6lNfNZepjSSrO4jrbh1t2dsWS/uefl6GPZAdqSSCfwGqYr8f+0qvJcyHbik
NzU9oHB5thQUyR0bKaiMwMBXa7yc5/04odNDgBEmgHPBZIYCpIbRBS/IZ9BGDSpzpDRTA67agMZF
zGlGDij97jOgM2FVozLVKW2bt6AeO2ypFHZi7W+ICkA08xkXPRWpsNFnTeSUJCHWS09jzwPmPKbq
jAT0ud1ziAkCNDYHM61QedAsKkkLO5tpI69qCKrO2PANllq9NprtAMY8QbCt++E5sARCOF30IBgJ
gnRGJ9GwxE83Gicjy15BNH36MufVRegtKadVRIH4/Rn6jHXosNCOwwThDUsC3Hwbkap0meIRZAas
uOWTJJ3fdkd3Ehhm5QdQQiQlQiBHK3Xi4HbqG8JofBhqjC3xnLXzeCpkFNhUP6LZC4qJ1OYzjkdE
qmMmClKvoa6eDNVowcv1NRshqN1b7RcryjLsp7zO1+l6jdwMWWDumP2f0MO9/oZfKH2ysIbXDBzb
d3uzJxZZumghWJOO8eluSP9Hl/68u+VqqmNypTrRp20dVYEKa2O9hc3Qbe8ThUR2XALW6BkWc9ui
SMQWb6Noaq3V4WQEoAR5FjbgSXCVar9nVflVSUT0mS2l4uEUb6Lqn7kMi7L9j9Tqt+tg0yV9HL5m
niVkvJTY7xxNXiZwQkFUZOFZzreEI4rQqeN+ivEpY27qpSPjRizz41kWEa5MmGc2baTxPGCga1GF
lL6VkDFmBocN76rXJWGnIieUHJG531ZQbd77nFL9E8sTek6AV51uITUqOHZICkb9/iXZ2O8IbI11
8kInoPwPN9dELsxl1lH48j4GA90FNLuOBvbcN8ajiOwrIeMAStelGpkHabPrapppehqrCMDJFktM
6uTiRyI964KKxlywW87OPyp4p65J4Uj2li+h6JzKBeI0AlKVPWXVTWSeQvnxOpqmzRIfI1OQPW/v
qTex5BjCiyFwaIMmUvLQVPoTob6hFMSL36ycMNz/IAeqfl2gQaKxywN8Cz3lMzkcxY8LUT/Vk67i
kJoEm7c1m0v1s5bx071fqjfrjHeXNhKDYjPSTPqSLDnF4ep9MGuPAaQ9CeopkFQKouRcp9TkBhBp
squSkAJ7cJWfZGw2wvCwoIBTzbexKBbgOeE7Cesg8sLzkeNtLYtPZ4iCoHNvN9o/Q8/81E8w8N0H
y9PBfV7ZTVs3UoiyPPVvG26hGC5B57Cc8GtrghRymVkwduPIYpvYcWfTvPMwta5OfHyzHqeQNzrP
nDoIKHMfBQlpZC155JN7cUw7len+r+NDWfBHrLJe7tqh+OxPsAwLmRTNdeyEnQIBBqQZvdkDynDR
FXOmVrrn8VfMv3a5awMQmEKv571RKKlKYnJqNe+XUuFq4V79cniNRcWSsGYstnM4C3YlGH0aX2Eg
OR63IBPjzrqE08PVTh8O869t/nsHtPvKelvS6UYnpyGz7w4+UYiiHmK1YybkQbXd89H4csMpWw5J
XILgf0wamD4mf1CWMmDvAf12z0i01puCwZMZKMuevcmHhWyftsH6LLGgAvYWQwmUo1BTmn329+ST
zPLksRPaY/sq5DEW+DsAhRbB1jOKNmIaOQ7lgO0yDbhloNmbqub0kUfvycQxJ6yXfKW4z09RFTEC
giUOlN/SXEiTg28N6dHbw61iXUKLN/7pUBuz5eGp1O1ciXOfnPQSXIlya74qN8Hxt8T8GIX+gc2t
VotEAkyj71GGwehOfVfNy4M/uwNo17e0Jz+EmRGvnxb5GDGtKN3ivOVg/rQghctRmmtHjSFj0k5C
w5L40boz8/y1zVvwZB+9mmPn4x8N6NjOp41KeVbjYgH37RcWti4SwiRKGHGA/+8mEmd1INgwomin
qqhE/uqf24XRMrYxUeiwRkthyfUpsiiD/SwZqzJzSJnX5ZZHbrzHmXJaukAh1YHcAF7v9rrCCwBl
fWaQsoObwfUYGJtd3V7Naf5EKP+SV51gM3fZxvffVVuXaVO3ZZktMfuVCsls7WdNKguHD1C7a7IN
fKfGwv4gguPCQB24kJidwHI/UGRUfnYBkSUU4F9QdER5PHVvPp8l50TYEW6wjMQHo9FoJF0IYw1J
+l/IGsxNCH8mGjQJDLSTk7zJMGDGa40ByAe+ldirzE3/Bg4GCB4x5Qh4CygGnDSXcG9JS/+BeYI0
pMkigJQCqXBFUA3i4Qd9PO5yKfhhoanqAWEWqE+TxxGlvByL6u1vmE3KhQyqIAGdMWjxnRbnpG/T
hRakyY5Gh3CU/FLMUsGUAD2BDCcphJConv4inU8zD6cs5pKS1nBRjcwEiweVD/4bzYECmKdALPTB
TzhF6V8S8Lo2PIvwAks9zIOgfmASuOw9t4e8gAx7bI7GPRX1EfXfQgXDxd1bi4ZRl+fx9fFKVoDq
rkHOX1kZww/SuERy8QAehLSeI0XgWNf75q0fA9XbOJVjDCVgXzpHutUU34caSd62J+yrRcq+w6wB
tks4LJHPTv3UTBTlSbz5DwBWmxP3AbyBh+LD3xoiT/UHfE93fM72qGBIsdXkRUvn9cj/CGporggC
1uQTE6Ycm6mhPQbFbUny/R2kihlCheWeHDtfgVniRyDG7rgbKJQjMQ3tCLMEvmLP5zXUoIixtwNG
qrVbuZMmxE5p0WdRuoa6xqtCTqbIi+3CG+frrKfA9yMofzq89ffHUTOk5GeGAAwVpwL9mlC1iZ7N
PnVv+YvYYVQEI+CxfH7GAKBy6eDw/hHViAcfawN+46l4u8n62mtVVQDBc4jqe8F3WqiIfuOlmNuz
/O4sdIsICnalwndhy4xO5FLtlxBs2WZuBMo3TwJEtktTMVKmDo5D5krBn3QrP6ksvehw9MepqyFq
lxpYw021LG+HJI1NLAcxKrPapnmKnNCxV/NUd5lWUiUWOs/g10PB1oiSlK6yUZugu64yhXshtkuy
FkOGkSSMI7cxRSqh+/pKdFG7xczoctF9oXtr9/o5tauqJ3HO7n8YfP3WOHTnRjO4lEZxH0BN8HZq
m7YRizos/mKNWPT9YsVEDau/fUQyABb8WvhQLLVtvj7gfr8LptCHzU+yj9OjO5dVK24wMwlDAR1Q
NNJx6muGhiUtcA18GuoYhO1QbJtMXzPjB+hBZmRhqX7hRmG+Dcwqbm4pFqk34UQF+pxw8OkomQNp
n+05OOR0/lxCMU+gJIsZaVaM43ZmoOBLFTBTj2AA4abngEjsreZ6Je3hni9mleO5p2Eb9S9jnI9d
2Plt9vF3sJrz11SU2mwYOKY6srQuMR6pzV0oXOFeV43NgLiqGWT3xgbcMif6zkqn1MhhUSuSbM11
zmYST//nQfdhN6JDsBgNZbj2z3gXvSbELwqDrCpgdkwZ4/qgTWqQv6hjWHBtEFF6+qxlHFr0812u
BHvkUan4a5Ne0jpg3nmJN53h4XnkKEd0GMJb6OYWUM9U++2uyMD26mM3t3TRjWJfBrVUUUHMe7O2
1wq/shKRA7Y3skS/uo9fq/GfkDg7WLUhfPZSjYluaKMYNEv4tdZqABz5fIR+XKp7WddVr2qt4tQw
+2vD7ma1zP7uqLTtHnpQe4DkFb9zsZkAQthJCAngfdAcmtBiY3rrXjV2U9RZo4bpuz1EI2OM2BGl
6ehAV0aV+1y0mxzotoZw4R3RgLu/KosECMUtCDUB4qU50KZgti0CH1wnALq5Fkd16ezL38FQuV/G
HK+9VyLGEOuuqXq8AMBr52k0MzQUqPjF9Moe28HKhgEZQR0Wk4BuqW0U51El3UazpQHRDUmCMCC7
E1Rrj71Qxl9OdCG15xoxtZgaMMnRzsi/Tf2xhocODBFVsDKel6KDXxjBS11J2FyzLQ8JhY03Jjcj
EvFm1CDCcv9/Mmt4PwCYbSakpGLVzPUlAwHGGKYUO22Xp/oY4BdGAsKhBx7rwHVc1TEtuCjVvyww
shkSnCcjKnGnrpXyc9b2HDskh+AyfJc1q6Nd6/hE8+m7JXrBK0xhu/R2nIDhWblGiU3HFDv0G8sE
65LiaJqdR9H1720JuWveStWm1xkwyVfqoUsm/d5a5dCzH+ca5SkkAvPwj803VptWCN39qvqmrN6r
Jpl7pivgulqQHQdJ1kFzYK19kVmH+A2NOkWcmiu3gVt3a5hcaP5ZkIfS2UXKsiOnEJvrOY6WWSu/
9Ms0cGefgqmz6Oh1qIgOf0+3maVkNFAZj1uUTZgTNtl+ToOKVndcI9P1P1q2d6fAS2NkFXouVn/y
NokXPFNisG5NJQ66MLpDcI2tnnLnnx3buWtB2Acz9kOhz8bCFkZJtIxzG8ExhIpIYyY2FOrcbJZj
XhwX1FQBkqrFq8k76dGk5WGJAAv34Jp2zFR8sPjica5wj8iNS6du1YYnQWyJnfxWexnNwccTF0GO
7M+rJPC2DN121Zp0kbPiqgW/HpKCA0m4qcqgz75qhJJBaseB697pwVgYK1yMooTSxG2KsbKQXxPE
FXJpOMuCK9naHodATsnnoUwcwkcGEr3jxSCIllj5W3jsVJpOLhwcw/w1oQpgTilxTz3uju0MQBGa
NJzmrz0rorVxQm5ISPO0zezlQtXL453p4y41IWITCl1Sbi6YigpvrCUJNAg1CDG24820FU3Dm/hn
tzkXPuihycqXiyh+ReRawNPMaCUvdDH5H3buoV6nmP24LRduO1N67DY7DBmxM0+P2EL00bXvhyFc
oaTkpabXHWIsgouMo3CNW2E1SziXhx32LRXYz7G04B10mR5Zlhn9QWOXZxm5XA9gSexR93eYrmVh
IO0G6R2nd9CaVBbRXFr6VK1M3QVNe7sjd/YP9HTK7H0fWIrwPIK6ds4wzzns3lr8/BBDXdVZzqAa
hc0eqjoc7dEe56JMtevWtlcNhJ32n2oW7pUOmroapWratllWm/mtLbMhdKKABif0iTIdOTUFgmN1
+K3IwR3132pMvGKfiRfZaACRHesdcPieBqhbRfwp3qclAK4v7jsRNDaHew+V8V3Uet+sU26X5U4O
k4E3QbVRpEkThLHOKMhIZzg6P/BlT4xehH/+k9WzEozTi6yk1ZnLLRAWt39ddgqAjjZKz0EhaTHm
ODCRGQkMBASQwdN1O4Iuk+M6+I+K1iexEddslsAconDDwbQ70QJReGuDNcsI3ymxzUaUGeJ3socH
bAiKDfVRLfYLVvvCO7uvh6s8lcmsbNo9GcF+mviuXnT61qRehTS0jLZid8nSlND26ZrNeifj6Dqy
WODMnI6qtWOx0mbI+QhAn+knkT1HMcQfC0Vqv2p0QOEVMYOMy+X1ffc5mLYLaM2P7TfnyqdRv5/G
Kehh7njJU+9fs2Z3exh/z8recEPDfsX0nNuqQ6ccAPppVnYG+1g0gWvRbEMeECOBjoCDwaBQsfpQ
IZ+R6UoetHVO/CTLwL48tvkAvR0qIk7ZRrFEV9cS/b8hwH5yHD0WKvehbX4f7CouTfF61HLbXEXp
/ZwqGc0U834gSHCG2eq82LW83DqECsPXBMAqNgOd1SSbSpCfxNQE+PuDEyeW6mow6j1ql3c0aNJW
Hc7NfrPN58IKGmgABYtR5l2QhocIoC1ixo2b4npTBq50/fSsnVfwKxr+6NHjzqK3xDTkdFLaIfLA
pV+FwjGfXdLAw9Fn7+gzRQ1cScYndmU8OvZdaxPw1bem2DRGFVJen/1WLxjYzZNOH6bt2rSQBycm
r2F+wDvBH4eQkXVHlQ0ckjgyvu7Rt3zXuCC4SOIH5MMq00vMbKGH+6l5HT9hFAtGao2BhPJlIBlO
CAch895h7cUbsalBSDU+54+RtGF8i7jBMVaDZD01iEJqAnDaexWEZ0jRh3MuF0dTkRgtwSrjRev8
xJGaTGMTJmSn8mL+uUfu7jJ+frs+jrRdSqX1CmEpC+usmnuTGedvehBEy0qJyoxj5NMVENsOxTvY
aK9DP3SOBbbGJIs2T3C4mqkbwXaKHHfcTLkX9cD4yh6Qm9gq1uDotiswbAToPwZujhnRQx+ClxwD
mQ+mKlM7LuykuBNppjXO7V0sK62F2+Th+aRjRc3WTQxtZrUEvYJW1lNdDlCTWng8R2ZB6TW9Lhvo
3v1rCFAdzYk4kkU1AKNvRcUIIbO6PIMvwMx3g8RJUhkqBeYqdKSsD/autAi3x+f5k6Gs7K7pxgnC
1OK2c+xeYKeRNgPNee0rV4fSb3aAkRCJtiNP+6IhiB2pFGZ7v9HGygluvvU0pdrWnO3CE4Kd+Iif
3rbtVB810tOdM3++QvWF8kU0Z7sU1T59MNxAPvOrG8seuDj+/VSn7NArNBN2l9qHYr5mRu8fr1qv
TA9SoGnmC99boGP4WZd1isPxYb1yYDjerLx+R+MB7nQa+ABp7xvBrpRSEApQ9Gpt+N+8JoxeaKKg
eAz91fn8IwVNa+azG7LccOENqYPmYdvWoKSYYfdDuIgeN6lzlfKELiZt60obbU5CsKTzVJ6mMTKy
o82x0BhNi862XJglJsM21i2NR2J62FIuljKr9Pe50i/4jgAwNuBNZ7mHuZDxMWBsp6VQtLL6IYiQ
94hekaL+NUUPCEggBtOtGyvlnkbcJO8PmmPnEe47MkeZh9kK5vqdP4UDAeQtUtKxbUYqGxYPQ8j4
I0Z+JAuM6pVUp2Iedwcqr/N8F5JY1XaubEGBNc7fFDJS9v7AHu8Cg+6IRHeJTFznH17eTZZ6keNY
mverqrtbqUPhxw4fgFyg44/+L41Ch6yko95Jp+Km6q11x8tu2S+JcdAWb7qwB+M4t0JeBPZu7ibD
vk19lcUwmk6b8Omd2vIrn9LNw7yM/WLqmlnrfs5JShFTTHCX9pM5jKAxqIScBuCM9aW+RPFWVWmG
HeVd9D0MZlayipGVhJqsee857wSEQN3XFQGl+e3ysAk0mb/eZvhuig2WMXTHZxZ42L1wv0autGv9
ruBxzwdn1FmZij/zX9zaZqDPWrx9Vkt8xWUwBNzgm8hEA7bVGrROInhfzkWXD8wSWAet2fN0Kl+C
Uett+mtuJYVIdipWTB/f2aBcPr450kqevnObaYG/GK21Eyc9OkBSTRCYyAPnglEnzcw1n4Jn6s8O
YTTHRCHKc/c1qYJeuOJobkRIUqce2sP00AgdLti5b3rqBbVkpNUNJY7dqBEE/eIJHsNXD39SqV0E
AXYJ0VPxIJ6mN54x8k3yb/aJESWm8UOorjkGEfNhfquRZmnPs3LNdFvCeeLokjTrzt7q4YPGHfdu
GlYoxhTBrNyQCctRuIt19/2wT9cJeluj/WItHAlmqaSyMKEPmKGKwgOw0S3ovjqhv/ourZOpGMuY
3KLDkp5IcnFvvLbW5+EmS1XV4U7KcsyQ9kAJ/dJ2wQjHqRkKISxYN/vwtdz1SSbsbOkkxcGqPtDK
4SZfyc0lCp3wf8S6PACtlZ8eQxfx8NyNKXggopCE6q+O7QxUToUMUxX4JCbOQbsxW+Za4XIcfG+U
UwvhPHEKyHEzJcha+fd+BxZNMlUGe8j7EsVPwUpKEbLOdDJ7uHpasUjYw1KyFIzDcnj0fQwAtSdH
YRW5LmJIDmvkUOQJDO2DHeut3Y36DjGOfBtLapUiiBjururZGavDkOmanKN/hA6daHCPgi8/dRO0
X97a/vw3Ho86ZzXXdl+cpycwz/SJeuHrXe/oqAht+0HBuI2oDdtN0X0rqw/y+lw6xhKCqJnIaiA2
kuF+YAgvT82Yparr7OAkbDGOQEKaLITeR2TRAmtpsTfjZH8xAtvuroZ2Y/w9Ryxs89Jz27oTvFg6
IWPegbhG6v88La1wYO7wjL253+ml55BV6MzzGVesgPM1U72LvxfpCy1PQEzFFvLkJI3RrDiBFr56
ooBCkHC0gPEcQLba664WpwYSEyazz8/mVs+Hs9OwjFMqVBXHL3HWPWYdLRAlAUo4pTJx6s9qZ7w9
f5mB6CDGz8dJGtcq1Bsy1/F4EwKlbARZkTwierWy+qFpm6mxwkGzsZ3NDsnKqYeaYJe3azYTMx/v
/lomjo/K5C64lkpPwu6fpt+n5q0lOcujRU3Mlv9XU4NdwrqJ9tHJI3dIZt2yMAQrx4uzhqyglobo
+y6j9I9JDwrs9N1TIFhToEwNwZ44VivDdwFC5YNQfkBNd4c+OcTxXOYCQoywYtnaFdHvNgo+qSXy
1GtB6vA1DPUDYLPtT6IIqTtslj+NrQ1aJyYLN/F8ibnTfawnoWiIuBvxi9Cgz6AUHNX5BsRwmWB4
dtMSKYDiW7ydXcqsz7gkUcpu6KmpcQunKJiTcHgOzmzxBIU4NJ0Yw9UMpstp9UpgDPS4yW8XM+U9
9c4qg9zJbKW9jDEJ1/Rfk5mRpl4Q/O36pvQ74kb2jeDz/w/yynjpOmh2Uf436fhhnzrMU4GPS+o8
CkTrEh2UjzAE1d+t/1NPOgpLWclEzvOXmMujO75hB8MXRTznDeHBSYacIaH/WV24nFHtck/1Vb2Z
m/DuS9l4apRFfFRH1Oh13nnua/Nxyv5+NXlVSZo7Ww+hCHO6aokJwUfeiJhxDJ56uD/Kp1s57Wkq
9PDXJ3lu6h88GG6iI2l9KHn9KFWmh2h7a1hsjGSzp+Ba6inJwFH2NL9W7fBb40dpYovWa/SShNej
RTFN27SsN+WOrb7eXak5KszujQV3fRfMx8SjwyXoaJ/R7PhFOVeDeqjwGIowp5+O95QuISR0ipyB
tTyvnf2J2tns2d1Tgn9gP3pSg1FMUb/rKRC+SspdRGNDcCnpxWLcdCx5y07xuwu4iIXytgxsgxIb
OxyTg6Euqj2095vlSqhfKePchOBLkm7msaB/+S3W/LAPRPTj9RJcbjzQ36a8eCkJERI98/o/SU9S
wdVxtKj0quks4X9RDtTZHlg79Jp9z8cfoEWjwrQeka9+XnNHP9AYLrI8pRYzAtxYZo/4Js+OJcbC
1PUbjMtVg+YtkhS5OjJBL9l95mWWn5QFCZydMM7XfEgHs0mseuPJ0Upa1eFEqvhHTmbRlG8WQ99S
vpv+kPdGjKodd0UfHIscQjFaOiJPOcEGTsHKysP+XuF8Ih5Tfk0vjrosdunMX73VzbNHZtvvbihH
z9jFPu4XXVNnYV4ok8VUWv4t75MWyHvP0Z5WD0qYteGF4KIMfjcG/qHD35+wYaAG6YGqnkl/hiKo
LxguQM/CHshT/9wlPbHTT0+V6bi7BV5XQH6gtJ6Zg3/HuOJMW/3y/S31hpd5rYDS+SfK9ITSfc53
Q97k//iosmWr2zVcHugaq+hrPt7YPWKpnZLelvwVYxWAKDYwINUz6L3N+j7BIu/+GarAWzbKf5jl
96DqzAqvmFc1QpBNWUBraJxRCCS8OBdZ3mwysIW/DMgwc8lx2xnvGc1P3lniXrQIvia/f7rl/YBs
TJEK3ih3QnAQIvKLAx84VveJis/x9bkPZQvZXDRdN9+saZlabdRDrCC4G5nt6a9+IANYM2m52cZ5
SjWTuNlVrLq14pjsscqU9u9SOKc5zNLdN0ANjL0xqO6NnnRSvOsXzmXB9Qp/GdnA0zOI4zgv93z7
HzBOaVoRQTk2GbI57c4nyP9smTr0Uh8yBRO/ng2NdrxUHrMdVIYCd5WxdYvCdcRLS5jmwfKAcPRO
qWR3ZJlIRHcaXxgWoGMscd0FFeTHzPy9nzPPCiRf2DlRXeoxnjYsQ5BwhBLEum6WxLlOKWiaIXqK
5F5M386BItZu+VSASfXlTYRaaqVLCaKjjyeMM50m9kOgVDi4rhGFrmew73QU0uqZscHwWwVwn8ND
Ih199DDmhcERsrKqv7eQ6GoRRJ3ubWnWYfaFYo6p9e4kGPuCOQOizXEbVv5CDr+JIZAid46uarWu
5jekkEUdPnIFRyfG1BfNydqcTz1WCezhW1wt24pUfE+OBWseBhrcQIBvtd+ipY4O71qGt8C2N3cY
Y6B7+fUQMSFk6IdIHlEEH2TtmxH/s/1NrvPdUcgOhSKEVExhxxC2DKlb70rLiT3/bHqeeWALdYPa
7JxojlkrgIEzsgzratUwiQegx2D+u9WKm64akNf4nQ0chcBuwt8B+VBA2UpANf6g/M8TIiQLolIT
vw7kGHd/Z/MJ6x87qaK3ca0bjlX7fAus0LpKHA07s5/TLGr5VZMnQBhVNWbL2bhta9UlraWa9lg/
0r4xPGzhq45skpAqexSuJpCq/WVahTBfV2IyQvjBJ6cnrbgaMzI2MXbFl67avH2u6jZodo0k51uu
+LoqxTaWxG6NSoIjYwMhUQwwMfRPakzJbGeKWHJItRcCjiab5ERbTuI0kuztBMcnTpyJfxUdnajW
LZ+/wlVYyS4peB8uOdigdzdG/8jahT+bEx3IjKCKoW5T5uhzYOhiXvmDwxwDBEwKG3c7o7V0OASF
8JCe9Ka6AlQozaafEjqgJ79U6fv49gRWdgL0BqIwiaz3h9TbfSipHyMDlaPukal/F7w2W6wPTw8B
NndBx7Z27vJajiMEQBo/Pxg6LIFZC157z49xGMm7qzA59W9+OHd/v1CFT3V/dgyCHHXoECKlOL/0
fVai/qJqnTrAe5obwaY/KTyxCs9G/NZsU2zDMEzhdM35FnseTdNzAfTER9dTMHk5SafMwqPXd/Sv
aSF74IaszVN9mEJZjaDcv4vwdPHfrZJg2b2UAknjj1iGgJ8Qb+CB6vawouZQZ5sQ1bjYxw4BZ2t0
68O8wNQhA6kuUv04+EUsunEu54xsjsmUO66RD8JxMNYrAWrd1i6kSWzEo67XKvILVufosL4v9vlP
MBOTFJIrVdaiWFbilF8XmyYno0VxEk3RzdKB2e34OO7hZGwh8zIwr8Y+zrRYOEhiqRyWucp8ODk9
9OGO9cTY7q23VMJEHVWJ1eFjtT2yzRDnOEqDwGizFCBnFr0SZlxI9VN8iUePAW7KNs9bQMTX26xY
3/3awDvxAKgo8PDhzekq4O6kloVY+V/CT92SKzdEv9Th8xvDg56b+WQe68XrN5QtwKNibCbxHIIr
Hjm8FLEa55W19tilbGdzGZO0bpDzN6t4uRIqcSb16cWQF8gx07b7e0PQsTE96pLiVCtMO4U9w9iS
N6gvvy+GlKgNP3W5wl2kXS0mQM1E9KlP/pS//LNommMcZYQ4GPhtpX+TbPFgbIQfpjFA6yskB1q2
eJFRdashM7Qirk12yG0GZdm5ZcHPdwbhOP7pACUauIIfKbD3ZmJdx/2QwN0XskuiskARIvGSvzSm
HNCnV/q+d95snS9AwjhMKAL6OB23mefak2vqScsVFbtbVj9a3vGJz4Ow8J76pmekjBrgjkPy/OEJ
p+xlNjbJSY7iW7TIoQBdLyMpUd9LBWHK1Xqy/BNxHaAHNenYekDB309YfYfaKU4nisiK6htJo+Pi
G7A7B4BcEPHhFuZArG20EFpKDf5Y/J08OEvfhTOb4FoB4Tj1ZAbxCBTTQoDgxWI7+Kxm64b8Lqjy
8229PVu56sTHPtqLG2+jvNpVtxb+3uIjBkTYGzcZj88/CT7zrZs/FNHo7VjFB2LaJimAOh672VLR
08Vy0ckd8JLBlQwpSLlAT8573bEIFraqeETsB/fG4TPZd0Sdq4tj4VtzxVMTj1IcnXGXEIx6m1ej
010tAnhVb8n0bCXSIehb+ESUcJkP0zQiO9oOUaSV2n9eiC/oo2rC0aaus9cCvXpCCse2W4Ntej+j
8pxVZqiaccG88ojHWVuZ4S4UExkQnG+4H9rc/WX8G4o8sQUu77WrtgtYuotTWj4GVurYz9zoSf7s
FBf5rBSY4zuRmkp+b/Ryej5yh37HmIYoe++W4r/rtNAS5N96cfPAsyeFJ8+Bd57nnSfuvMeuaVYq
8ZSkPjzucjmIm4LvAu7EB1fTjyzylDkS//2p+ykuWp4/VH85nRWmhV1HC/ZBZnPIY2oI3w3xq1KQ
tzTylWfTstufPDExJLt//GQrDIs9UyQoTS/c7NEMg7NlXQMoF9DSHNbMKwyv9VPzxAxTXo8MIbON
7dPKDI3QkxaQbON9YrC3ll6Z9N7oqHFgMftpnTNplQ0kUcauTC8U99FZeSz8Gn10P4R0tgErLLkz
ySHgK0Vw0HLtIUBf2/he7vjygyOtDginRctUFz/gDXgT4b6OcCm2p/cp8gJDuaYpaouqFud0hVrL
CIn5PrkTHD2gxfsyxYNAOjxzgC1kRTdEc52ld+G2dyvo9Z4aLNUFLP+Rj5gpDWMVAwiVEPT+2pLh
vTPEPCBSmHz8HMKZZgyGOA3EErh6DWDelAH3NTzEoohCilk09vfXhECR3taWb0hvfHos3794EmU1
/jBtWj4NwflnyWAPzhLe8xHpU4eFw//QX2iXpPcHbIMqqcKFOTq8MH19O0PhL/+euAUbLpx205Mn
NaZ4iNlWZEgTvJAPzw0sTRIh1Ssbt9XV66CfVEDt/rm2wtgObVXfIKrfPD2lzotSFOgvVdBtWFiy
5HBE6voBcnGqJnrdcCtDkeSkVUMtbwMqosn1fWoqVO7Em4hZXNdUj6Szq48Rmjxod5hcbFXprYj+
p0ZhyGtLTl8bB9ZNvaZ1rtP6AMVVw7jGKcZcpbSbGrOLNBtz5pR6ipseclkTnMoUGEXLKQpLVibh
eomgY12vFXpmF12IGnNVCnCuyb55Xfl6j9+FmrYGMyaoEmPeFBZpwvwBBL5i27Ld//FzB6b3Sc3j
TYQJ42mgNcMvyT6m7n3gvFD+pvv4LTYLQKx0qmybG/S0WR5Bo8lIqXvTrrDlFkb/OYPYc1/REB3V
l+VSdsNaiJoLsAN2dGPkMTU/H87+KTRCqNxz61tP7M2v5JPZikygGl1LG+XInw+wqYyQ8YDkPanS
mjX9ScQiAVnnrCtL/sOyeHYN6iRJNJO6jpiIsK1zSWpAt4JRsaQ+xU13/1Y7mhYgr5lfzLIOwsx/
YQQk/Dtr2RYBMY7t/14kwoelRBBcW+JCEztWk3RxxbkJ8hyAUBYILCeYCxjw9938aHCkOqZZuxJV
c+3zA2fZHlRIeOcJ4j8AdqsB1zxOg9u68Dyd03MWWfGzmQZo/ZZObkT97JSyu8NQ+/4by1Xb8Xi4
mgwHEOPOCXzCMPVrhwpSaeRDQlgdtW/Zx/did50sq/3JJpxK4RPP9M7Yzlfc2hDjKl1Bk2P2If1+
zP6XfoQ79t8oqHI0bn3gaNH8Lu1rCzygnMuay7r6ZKGbrwMRC6s2TMcJGK7pNDoxsa8bD/0ICx8D
wXY8EO/thefTLi+IMsTDuMUMch3vohSvmO8YDBBT6pmN+j5m4EekNQMpoF05BK0Kou9w+sP6AyuO
m+tiGRnGlNjFMtVqPQNiFYAa/TSPFNFxBslkuQp5Dfs4atc5M3/fHuZ79bnnrXGI7lZHdc0ez+nw
SNCy46X2k5pnmG8ZBYNyHVZvNRPTMB8l6u5sBrxi4XnnsQadepFq0veLF25MDR/sP4guJugcbAJb
0qqhB1ZQrdkJ+Bw4oEGtu+aRUSVT4oyCk4GnEyXLo1fYrKkWVRund7yVc6yEDXRiLst3bFkYcWVy
7fe9QYhuF4jkMetiQPp9kYBkcy20lXxR8YKtV6R6hRRuxc9cR7BdTj6SJnG9OO1H51RBDI3uT1m+
qAn0ECPxzikGusHDizHI0ccEl2uyV6w9W0z7q4TVZ1PJes80BQ4uiz+ioOGcKUAxnc3iazdm0OQx
9V0spxy10Khg+TkonL+mDlmpVJMJC0Juyomv6mll0F2IcRoQONB3gC2j2v9x8RCgj6ZW6PD9XkBP
7Af1idGj2QvdD7Q/olzZZ/XgLbNWL3oAqQJalo56AwzjIoPejNMsjV8CuUAtFw1KOuqMyzY3Shsx
D8eh6KgJABn4jq8DiNJ6P7i9tR4kR59JR8Hx6kZ58l3e0UREF6MuHgUK06CjGS21SC1vLZr5CRb4
r9t39KKMOrPMroAqaLDqnS6fGUlPG45YaaIop8n61nsfl1wvrr8X+je1h5YjxmkTVVOG/RQpdd04
xXcqrTkpzKZJesxJBqWFWQHiDkoXel9WDrca6km3wlQkApk8fbTWNfThhqX7H0lNnAg6rTUz5FQB
HACG9SZds/jl+Jy825cZHp0GpZ9OCmMrIkGcE3utMAf8vAP8KOkKnu57Hyx77OJtZ/8yCvr2vsHj
70s21XD26TMxeQ1jfodxb8ctA3gGjrJp1Tx4fI+r54aZRWfI5n7XRlfM9VRxLY50PJUUj6KAHbiN
i98NffITgq5aBNN8Xgo1kPj+DhgbgqW5ma6FxKhMQw9/cNNhxG8udBSfvWq7E7ZtndRc4uMO3I5+
rLPhfl8CljHCrLJrAMmX7UlufXGCGv+i3/TpbN/NGVA890IXj5f2wPRXVm4oV/oU0v1XT5Z75BZH
1vD9dFGzRxo4R7rUMEzG/WsfNSS6aNeJ2QXHLiMUnv7SD48YYMlgIwjuL9bBAn9KMmZQHP+T2dU8
9rQ3nsZlDe+gO68PuIhUklnTqja6bRHan1uAvQflfBNwFMs5gn91hthz9XqIY/SxdRG1cjhxjKbs
yGF08m9878xDQHBDIFYuPSsjdKjggLYjJk4hCiinEMioMPeyfxcjrxxI+h9z8kaucnUviaGY4vvF
cuxOSqGv+OYzWgcGuVRkzDknYTuo74KIKUhvxVMgWu0CgnStJ2wG4iUqDEJ9WQX3brpUS7JPtEnZ
CCCyMIHdZehjj5zxU31WhiPdNP5/rJ1NO0zCu53w8DAMiCIcRZeGdK9kx4+NDoQgjn9ViVatV76J
m0d8XDY/v0WEmLVVYwX1uHTBOOyUL/5XeydrqfIriBXh25ZsKDRvkYfwAE9rOtd3aV+pX8Gr3CKJ
AnVexobNylg4C2Ozg0HVMevVXPOoVfpR/6zQDKY2Qs0jAd40oed3lObr2j3MBDaJnZMIfj+b0YGH
mFi4txuO9uFW/GwBKfYwpAm2fK3BlrNKuaV8rsA2i6TQdklix68JGzp3q+9moPQrx4GBU3Hw+1zL
El133Liu7Rwkb6syMdWPmAh3CBv2mncCgNl1JQ9hWw3WRpDCHjqRV2fCYFow2pTpO8jNWxnr5lTS
lGPgYsD40rtJ4g8Do9S/6Tpjt9oxQzsW5dHgVVMtL9xxukyInfQPTSdQL3xle6kVKTaPj7/WxglD
usMYSbMbRKZLiAjs158snKnrfiajlFPaytJcSMlSlRtXggTmK5UGamk7vXQzke9wq+Alw5CCFDws
8Pa6CjPFddanzYMZrYqrC/O7aPtWCv+yqadxAJz9BqJdksbBGYhO4h9x+EuWdelRxq7ewHtyN0yc
h9bVGdtilxWf9vQ4vmm2EQGt/+OrgE6573YGaTDqp98U5YHDmr24dvbXf83x288LtKWXXXPoeN6D
hUVGx0K9XqNaZvDDZ9Jvnf6euYq8R+oeLjl1n3rjcnJblnQEonhGqZDH4PCS90H+Rz5G63K0+I7m
TDz5dOh0Hbrw+XVbQPkn8XT+kLFBMUF4xN80Bd53sprfSu2ETbuclMHZBnjlZYWw5Bt161LOqdKS
5aUaxsHTY4iLdAWCjsftOG8rpZI8L6WygLgThmY97sR983vucga+rcYQzOu1AVxkc75eEyn1RuQi
8zEXq5xsryar2WL6i4LFk+2bSw1nOZ4RjNLHjdfgABhf39auZPXFhS4IvTU00FaIf4nyDYaHCDxy
hnas9J2d3ZfCIzWGfP8rrn9Uo5dczkfOiNWPwCu1fVBl0yaCR5yqbsZTTAGlyEknQhRmPvqd4ncD
mwRu4anokx+SnYgiRSQC9GgQ01JhA3L4eZ9Yh24e8rMJQ4LCv2sfTzcObZ7bhY0DsABqlrMqpB2o
Ivg38rL7OiNwkX8FXC/cgtkFoXPxGyZDktfGMvTELbsMIPBStL3oDQzn/a+xktcsi0GKjQSsZ1cl
XVy01nCHsLZ94SWCESGzXLRbg83kp8ql3gkHI5sOhp+qalWiC/aNEjSvlDxircgFb22yHVIU9i+x
LnBtvuWe8YE8SU2CvkoeAoXIVEEeVfhYIH3OZI3MmIGtOw+EU6exINCLsFnSvG57ugDBxk+QBIWa
St29pVgaKbJsL5QAllfvxjnJZPxH4Xh6/0db16nGfh6APLI9S+/f+KU30ndNvCRg3VvHx2LVMAEn
dLrjnhFgjro+BpthmMytVMgJjuUy9GGKD4EjNWHR97ef+YbywaVkwUaD702rTdnNPc7OoQqdQzz1
P5zDHJI1mqhU8MgE83SSY/XwBL94EB5mGV7Sd0Q0QPjWjMvhKVC4BTbKqBqAWyrkTv/M1u8Nbya5
gbAzcAXW6NoXLX5f4WEWdxj//qrpKYwt+8tUDrJLBRzARmBGVrHDGLthg0a5xBh6G0i6oztoRj62
ZcdIxazje0VDu0jmFEtZrMGJF/RBaUH4QhCMgmnx9XZYTncwrTctTEJj/ezNZ4r5NgJ3j7jSxjob
EgrClPoCwIyTZchBo/glmv2ot6XWG1vwX8Hvk3Y+gztHaoBO4bS6FSiYUsZQj3V5MZi/T4co/tpU
nkExo7nosEWazRUwn/EUarlT0qQS6wYr6C3xkwO1LFXmsW9tXz1S/wMZv3zIzUDsqgKDDzH32MJo
QZHNQc/mNZOc+RSVW6XsWilQKlmmZs4m93gY8ssIvliaPh2w4DSKV4Lha2Q1JnUvB7Md8iKENBms
7eJEtGwHJfEeKM6pr+eKGizgWQW5zOUuPeHxHP1UPYCNPPOPn+80B//PXixrNU6mhmyew5mA5IjS
FZGA6TwJ4g3X7qDixwVE5N5gt2tWnx7SnXZ9IlLjNOpOpaqcyvtEzEAbGbf1Vl+x2JnEPwxcha4q
4YAzKU7Sk5aGKNQfpdlaHjdTbqJ6j81Wy0vfXj9XRI/J/zVk++cVHg7JYe8gzWie613mRKjoLXab
3MUhKfbbrLIeyylH67WD9x/pkDDWtlkdv+8ouKfgyEGEgOPtdc0q/5S87456Ctn/ppYtDFUbHYEE
zYyh4mDwdfqTNozBBG7wch3vKCwNZI5rddWc+wEGZPcazp15/t9RkJPTG7PNwLCD60xi3F5AD8hJ
kUMghAtBxFxZ5kPeF4xDy+2MSeAr4+zk02LhIj3+SnbCdLIMo8+UOlrmR3yCom80g7pxo1y/U+7T
no2RPaw8fNcJ+CaEA+qXzeCQqqoKwVKp64brZVXE3aavVvdIdtkAPxRq0/0f4V6qCns1pWLE8zFz
WjnjsrXnJN4LZiB/RmZ0qeZpfA7TQAK9RHve0439I/ar3jgmOw3sFxq8EdGZbwE1v8PmpqSjD8Za
NvqnsgM0t8xbg06QijnAf06ysn0e8403zxWGA9rYDLHt00UrQBlcF6urt0ruKMrand5tH79tA5M9
qqdkzG76Inn2j1dn9XHgRkqRklRnCJBQet/8ayzJ/Lf2JrNWuU0h15nipTmAT1h4ab6ir8zbUDo9
WMKItBFNSpJAvLIsDej5HRYILsrjEZ4kCNcOEZRmfAQSpV++rJbdZSvUPKWCkmiWd2dDA/SpeUrC
NWFOIdh/YTML4mir0l94Gb7EVQ7qB8by8Ql/Nblzn1qlPHYAD84nHvkEkxC49VGybJnouAIT/2AN
bo2kWXemP/2Ua/1c8A+nVGu6wLl4XGCzhvI+VQdiMtDmbfwwNL1+xrDLr2yntU+e8G2UxJGt3iQq
RMbvBQzTea7/cQfNT5ytIIultqhB/L6oVKwR8PN49jW4D6o8h2xV68dznfUGxlygjHs3NU8e5mLE
JQGkJRdfX3bDFBQ9ryeD4qMjPSf6bsWHyWBndBVMutlQfsB4+E7jK3bGvRFe8N4MLlkneFy+b+pL
SqCVLbKrzhquPCgOr+2q7p8092/1Wcxzs0RGDq5t9EnalbvwkAYCUEq3XNRqUsBtF7QIQdtvz2dP
l5da/KYiUw72cybJyliwJRcFjCyNj3MxHW9mX9i/51Wuz7rdBgLD0Rh+iuIDCleli7a2/1etKLcs
tHb+r62vMkVUoBzRVJhiH40WQDo662jMjn0B7Gn+tCDxT0i4THmS4bbRULEhwM9WzCYTPGIHJc2R
KDGtCeeHqoOQg9cOS4f5+I5Hlqpz/XQCaFwpCkwMXCsYhLBd3tN7gq/y8wTL+o33TomWfoCRmhRs
w6mjG6nPi3eJgXY+YY4fzcXtkPuX/r6vIcJjS19MeuEX8SobGeP/A9UyvtuWWh79v4QxfoZ76Hu8
aYXLvN291BFyXS42BdVxhkpWt874pMvE5baKH9Ko7yjaQKCPC7BI/Wg3PnJX4d6EP7hoB98idT3T
ny+tgdVTcwG61BlxW0J6L0he2TI9y92yGleVhbhcmNdyk05NX2VD+xVqPjyf1PXgHw9bwNMx74xe
2nckVCLPB6zbV4rtEdCA7EhaCUAh30+57embscB69PPlC6+sNpJtkMXtHvbdvX8h2gJtm1vg4qel
w8t6TKXFWhXAVhJpMNgq0Msz6rvD0xjSub8152V8EFHh8NIp1AKK6VX/AQO11hiY9JNHgHDvUf9x
f5sUXkXhUCksN0t6eDdoVj6rntVgUAUNAxnxWQJKpKAKdD/YuDRCQT/yZXN5FB2su9O/9B0z6eZt
Q++F3S3F+3ELLIInqz3zBhQqiaVgRIJ6J2MxRXq8blSQqLK68K+jlT/2Uf6yeR59DAV9Z9Hn2Fr4
IOSIWMec2hUVlGWKbNrJ/84b9rKaMyRr2zpQVMlZ+s7vy3fKUsOt5xHVIfmq80+zi6yqN0Ni2zuw
KsIjsr8ufclCdaDc9ABZ8H0vNDZE9G0JmUnd0O6yK8w60cPeTbxTsnKobRggvp5IcM8GmIvc9l44
Who4nJFxwyVxp1MPImgdLiqOtbADrcC20PMGouqd8IZ0WpDzIpd1w6dFwi7XtgIdMRNtXDAjWMk/
kXpd9J/gfy9gP9N3w0rzUeWL7jb+BJQp2tCBOv4hKHKJkR1zZ+iFKgJiyoRJgOueqfCZHMC6FtcL
+zkdWmN/4J8dCmt09vO8lgMz3pD18TbEPQnBU/Yu95aMHviDsIgzplmboPCdUwjaByKwZMYm+0xH
8wASDGCBhy6N6COHNm0HjUroaVP45STlSlGa4f8TbRb2dFyhcAnmyZAGRJoGn+m6USPb/cieTDoy
Qa184t0+ewszBj5H4bDY1I9gMzDVpDuapZr74ArxM2pHN7d15o5jdJAqNaCti55NYwhpfbzWAIKI
pHEFXD7wkcbTUbKrqBf0WMcqyyjDSRfhsnyeFidCZaoGcUMlQxzt2bhStuDsjMrFtzfsxeRwzUgR
ucjN+lZH24MTjBREsTLW/aGjV/i2Hhn3ESvvZhW7Y8XRb1kDUpO720u+LmS3uxz33mTRY8M/M+6R
JrcVGqsbKkES9nf8YZn9YHRXY44s9tI5cKLWfqimaqGtkntMy/tFnWYZF7oxdVh8ymI9Gxp/mJ7x
aU5VEo+SYHj6m9/SApMvzyG8PkwtadxWCFHxyxgwG7kwx7K4NXjLTRLRh66xPwYey0J7xjf6ApgF
IGG08oWTRs7mu62cVtdtSW3c/qGfW7yTF9+wRVYwHVg7ermuFcDFxiYpNKPjijb8Ok6my6xEuNuU
HscVQ+OooAXOAUa2Buaxhin7jDr7M+ktMlTv7lq7QNJL6DvrdfOnBOtqDDM7sn8SIY3f8g7wtNtz
5YdS4Yz5U8f3RaHFZ792FDd3hbhfg6QOQYMWsTj/1lpy3aM6tn2EIn3yeXqe/PpuB6ua6K9KrI7J
cUH1fWeTH7ddAkqNeg/haxqDzgC7olMcj8S0dCf1CRBtnRv+D3knwNcEyDU0UJaX/2Xno5PvFf//
tGKIXwrzERx/nGvYJgl2jJyy358xWUyWgtOriIdK2vypzSAuCYhRBJYLPouP2hxinG8HbmJirabw
GMNElPHKPvNv88QbuO1jy0zD596jvEpxvcC+T4pYB5Cmd9BrQtUQVseV8ILWqr9fUXXmpgGmYg/2
LQNGQsTALTlkmQYZ5AXKUwrWCQudEv1v9l6FiSyz4idXnqVDcoPoPg494kKn/EPzbI7Mq6kvDNZG
hpxV3WwXJotJvYxW2agzPojKr2IPht2zjMUYTSjLQ5r/Xa6qdGdwFKXOv6NR5uJxuu7KCW/ipjw7
5uELTRalunAgzxWxPonFkVLWfE0jJBZwX5njgQb3bl9PFRht/tRXf2tJ0aVnmjqT+ZLZxqL/ECHO
Lc3w3Dltdsc6B8k12MjppgtolMqAtQ53omswOmDt/8oBQ/oTKecNtxMh1k6gEU0dRFp8+RUhiV8m
UYxJtOTGzeFymAcV3p/bc9oYoZIFBemi93qiTPgvIRrj8PHC8TkROMksKn7bGRTjWHMGskhlilFI
pso8zG0CrQPN3QQMYdiRZnJ4Id1/xxDpIsOgrOfRDedkluhPacL7K92pXD6hW+qQb25ZSJLWAtZV
OKW6cIr0NvAFbmRQUgvcLx1hT+lfE4lIdWh/YFud4hRurptY4K3ibIhjMBtQkIbkV+BZDUegUbWh
ux3Ocz09L3cclQA4T3h8nyOpUvlXKjrCKyhwcdMlFv080zduNyA2NhsKV/vEPAPAfya0wmzvb2+Z
Tvjzo+Y85OZUr785Uxs/D4WCXbI6rNbDH9G978vpmuGf9W0MgDkHcoRzNWlpqdQgWtj3KSO884yC
Yh+EVYQUv/PiundRHnPV2Xm3rvSxEdoIjQCNPOC+2+AMIicGL/nBDdmqeiLkuCId41RK1UpNb4zA
9ZrbqD33H598x8sID2PnscZwHvVNA6ujq3rAp7YHjuFNAQt9yWPujxfbqYlMqbEZElY0zXoJIf1y
DMP8Ou+8RFvZW0HSmduYO0/ahWyiYIYWcwUy8w8BuTsRB+iB4U5PrYqLowfglMCr8fEBhHOMhUlb
w6bJGwHWMqNdM2J3477Y5VrD9XKSWafhHnGUSWbdmovcmkZtAnWdQTp8lfn4La6gk03ISskt8FYY
rJBoswOIZSb0ApOFh1qIiOEgQDxKTDFG6UXrUM4pTTk77JQU1b2+ohA+AAP0X+RoiOT8LFZAVcXq
WNlxxgfVMENcSMhEzLgb1/od2o63Ie3h5V3RtTDANZFqKPDKtNresmgOIVHcbmG/Z58caQX4U6zv
pOYzirRXHicNhTG0r5YAG+IBBDv5hgwaNBnuC0/aJqszVqr8huvh0EsnhrNOp7EcYoVv1ng3Z5cH
LvrR44e80ETOboKe19ihQyQKNiDa7DGl6pJK3F7Cv+pvNmWokAedvJTp7PL/0DLo0ifHuBVsN3tL
wfffUaDEQkle9xlAoQ5jVtDN1uzbkZbFZYo0mS/K5PtcHHtfqk3sfR9Q0m8YwKlDDKDd7HHShVUT
mPTrIeLzmyaVzu0qEr3mZQGbQak5qlcBDtMT1M6+rAlH/A0KIjcAwOHtZ8UQbehaI7RDtH1JRl9o
Oi0aXkXmNX32sseYsASwiKg+mzPdsjbsgLjL9SojZFxWWRugMSIBhJYMDiYcfXREm6m4rGdlWUAm
LWO53hu9Oa5ETdwzCe6LRb2x4qzUcjfQ+q2xbfTtucXXie96bCf/kXkqY7SgS1SW1BBHjrGylTko
/t56s+aBvYkpe+RIOteEksxcIeTelgP1cWXwJAM233uWvXoBhIpU/V4VKVpu1pYihdgkzTsT7TfM
dmXxjnV4b8cSBWAKGDFyvZTVhfFC/x8Na55bznJD1gkxIz/AApzaXNVw4tQtf/42lIUSPnem6xC4
LipnkYpxI+b9sOu5VoU79qdatZ3VKWV86oqo8kUtCnpjGpIrKmkRhY58Vim4SPLCf8ZwXSGPPTPP
6HUs9+ZhCa65pXNHsdGGc4aPVsSjswW11YY8RufnAp43jlQTZdZTI2bHZ/HX9SCxWx94ubRshfau
RFCb/DPTU95EJ1/wavprjuKPnVQvZbiyBaKtodVvjTD1C5u4k01WKVkPS4GONZypu25lIqkSfpCC
n6jKaUQz/7I2QtPbb6NCEDeJ+S15lejgEmZ2k/D4ugUeEzEIkD/lLmkdMtHTFIVXZmERLx2wunTz
0v2zwPzAFdI7oRbmpWalTWBVEBVLBCftJ2sqBPenCudqX8Kxy2EFnLTE+81FMFIm7bQyfkZ94T19
JAUbdxcVF/eO3J7jzl8GLAgrQmR/wC0SIbzYRrqHRijh/8JXPKapPAMIgUbTdGuxlBwdDaTpvMBE
SEDIxhNWD3UJbQ9FDUHRRNuwD0AoInaWkPrRqoaqUZ2CR6DdatjzaUyeorekSu51Npkd5UTiESPV
j1L143efxiU3iNhNWAYvsiwOMrIcVFa1a//L/gflnxRNtxMxN2s1+M9by19PoCvFF52oG3WQdceQ
ASqdoQLaa+9/Okcc00o7XR3EMZ2tJu8wGmXkP06D6Z5Hize+rNiXNz19Yb7LLY1Co3vq04ZPTxbI
uCZKfslyYHwlGimJbyTRq7mywfCFLNokD6jAuSnYP+mduyLMPL8NeedMl+X05qajAVwUdIbv3Un7
oMd1wywUXhVTdBZFSr1gQs9Em11Pk83OldSZ0bhb1q2QVtpTXm0Bv1nL9+YuEmvI1YTil1re+IVs
DMhF6z7hgk5g/29ApWf5/NOMFfe1STCeYthgBVNryaOYSS0NHdb/K+xrgJa/dXjT91z31MrpIalM
QXHC65eAyFW+cWSBNH550bcP1TWAWx4m8Q8madeIELe90lDvAL2oYZI9yAvZ0Ubpi6HqlJ160Fxe
na/272uovsdroBSfG0nUXCq63zRufGNzIssOX4eL+Vs1q+EUNVEnY+q0Z/RPHQnxxlZ0l2VWELyz
1Khb+/okjhhRXG4Z7YqiYf+lfNjZoT9ZRHwdtd8UBSXAlEJzwvLRyeiDPPSkNpXOh8cnG0oNorhG
fDQ8hWkkxN3X80L9T7hMfc8df1BeFzqv7vIK4i+buntDdmbe9IJP8kpzRPh4S5yzpsPk6dU83Baq
Zkgi4hOGL4T0But1xoSjHCc45kxWM4t+muC3xxihMTkw6zEUqmQSEKjvHwte+ArFCB9bgZ8Op1hf
Pi9FOabZymeIStQb35kLa7GKmW4I6QNiTGFNlDwxuHtqR5/YRaUbdwcsbxR56fxdp2ZPuGPDGw5m
pgi0CwZUuWBS7mhX3Ar2NUqBF8Ran/AfSoia6ww0vPc83hY/hNgVxnV+PAQyJHsqbcQwpvE5KCW3
t8ChSd4rD2fiimVKRZRNM8NImObGJR5UPDxAnnPOkVCiwJJdzdQ5Tyl55yVy0AZE8wVwM0Vx/Vmx
2/0A9ip7JQANeHmtEz+adGRcGsSf6ikt5rIsa1sakByFW3lhSARmiVD6BiYbUzb0fYWQI1sVYTO6
6LmAShFq+gzDyZO5LpIjGUXBW2VrbW4H5Pf+5eElPneXf0gWY9b4a30/CoCYbvtZsyetWLx7gz1E
Ww/Nb2GmoOW88hYeX3/TgUdIRpVZEaHobKUbvVoHbgryO/WqLByQOvjS8ZcqNVww8WbnfXhURmK0
UaLaX1YlJPaVMz6G3+F5r1hZwtutXe93B4+T1x0vFDGzBXFjXIgzUzfsR6T7yAYmvZZiqHueyTHc
Q3G2LMIcCWeEWE4Qfi+SNaQ0Xe5THaH7ELszwHv7uR5eAbH5jaWhoYtUMqEm1+tpruaoVvgnWSiM
pr3u0MLf8Y/gkrq6aAjiTvY/2SovJTDhQwKWf6iTKHNjpd5jUCWSQK7tqxTHEv3IOFv/0g2C3XvO
7lZBfwFdDK1cViMmINEKBHIkRTf9VkZVWFfD8f2tzvPa/q0D5NPhJ5ckx+TBvSw0mT66VbH+CQD7
smii7XmDde5wNwYHa8VdW/Av8ALWGawjKoq1QTgoMp3mSspuGuk7kvFlhagtHPm7FEvziF+yQYZa
sLFAnbyX5BHDQyGdTk3D4qR2euWUcQgRt/YRyp3jeGXE1B92JS4fGJDjL9S0uki3CuzicYMsdKa0
HacsePFpbz+/nqarq2dPJRNYuxIs2OWTVCvCzwb07WAoLmlWlI8Q9XvMQI8M/YubuTu7KcAhF9bl
gad+fVU9UVEyE17pwnFMiyzLNU/QJ1al93MDNpcvxacVwRXevZANqEVcAVnx8K4Ur6wWQrQLij3z
mDz/kerxlXPY77wgqFppXeMjLjD5YtMZJNrEyGO/KptErais+s/u+03mZ/8rjmmKBDIQB7vYzV6m
5DzL4u7NfL+vJgPdefPT6G7qiYmDHbbDCZoPl/SYel8b3vM73gkg8ciWWt3I67dUpMGfCmApyljT
6Tvzk6FntKQ5deu6rXhsUrkDY5hke1SQT8ykgnBz/9wCVjv+23uJXdvBVQ4FeoJZPc009rcJNSI1
DHXwNMxPYmJ1KQu8j5WUHiKO+iZta5eMf2XA9bqJoFPRxbh43c8GhwTbiBEckwnpJEM+yQE7hi1S
yXnB/UW82TjmEq9+r+/IULMNll49Ptr/oa8ei21Q9+fgC/QxXCAVMeXAt/pH4KDmaor7FPjPmKyN
qb7qNtr52QP6y8KyjsAZpKZurcIzbEf7JRqZIF0qIRRSLQ6U+T5KBPSXK1Jfrnugu4dKQuQqYnS5
CQ6mS+2wFz802xZs/xKIPVI/3M5f/kpJ9B1tOpMZk4Amtf2+BTKC9UkY+Y12hFHYv4N/m+8jQPr+
xm1hoNqtm5unZkZ0ESVoAq2qTFcPGVAl5H99EJbsNL+rgZxSsShks7jqjNyWemuFy3YhfTyhgRbP
WGjN64T3/FH2TSgZpxC1oNhCILP1RhuKq8jVVLQtFgtc9swEZ0K1ioEhnYz463loncVvwbmMiJVA
cigvykTapochwxWRjDWP30uOGcq/jelOiVHmzr8x9LdR+5RWB9Yu152tzs12rvyxPoAkqngCGSfX
HKkg6zVHzz1DnpLtTux2nqkUoxYflsfhQt1Lg+BsEPNvnh4XWxhyRGMRqXvaCfKp2y6V61aoGAux
SPxCKSvUVFGOCjmPrECjt+YINvT3RqNK97e33eB7d7sRDKGNDYtpk+4ld2rQ63aysfnbD40TDeSN
I6KnAAavZJDJfC4EIeAi5ENawrYcqwo5x/8a/rzFDjXiP8nEDIkW13DIaK3XFvVzcwqZoLYoKYrV
9mh0TWuw29QL5ErkI3QnuFSuix3hXJVhomYQT8R55CnehOWAkZnP1b3dONPwvbHCmJm2WxCeeIpv
Ukf+wK2CHQtDwoM/JpysJjnRxpYZuOPaUGL2CnNp56JW+2bwNh0r4FCqCfibJdbbdLC+It86PpbU
pOE0sAotZJ4egzY0gYlesrupROdCRz8qs3zGILfVfh741Zui9JWG4BRgxL/QhyiHQDkl67+D4qHb
FNc87yH0DXLzDuCX1Eg7jwuTZy9bTZhXtJphFpSHsvgV5Bv4nBJO54w5qS2Kq5ygBcMg1F+kwYZn
T+65R162QsWSxtbCWvTuK56mB0/kfEJMzkhFxhRXXte/NMYg1nZFr/9rBoUKeCz9ycIbsIMwaDVC
lop0L76R95GxAueek18+CEv48qiAgcVrQQGs8y229mXm47Q8CRGxOpZSOpV8/1q+xW8X1IWu/Zn+
5NoOz8IrLETNGYrEH8J2tWcMkKNGn8uAReE+a3aqVFEh6WriEsX7WPx/LDbfhozeIL2fJtqjVtxw
CG+AEJNHXCaY7AxeF8pNEDJ8T2uVzuYBnUvs5KYj+n4nSnNPojCIpmPr4m0yurGSk9tpqJ7QVYLl
ZgWS15lIMEnu3igF5BiRa2RsqYULSOFElyNb+JBGqAsdhN6avV9zIKKgmr8RI52WG6i+9UaZNS1n
j/E+oRCv7YXPLQWjOnktCqMWaAAjDbqvtfXv5fMOmA4V
`protect end_protected
