// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UNnpa9gtVaT4aRyjPlxqLuJWbEruwicOUH2asFHN0eY8YeIPeT/rHh+vnPgJccKBPp/3fKSEocQX
6SLJ/Ih2fzbkvPYzh5i7oTE2iUKI08mi0KDUuEeO9kxRO1Q7krohuJuMk1bm67WttsGIGHj3pcte
EqE1LeDUtBMdXyVSzur7S0UeQFESSG9R0CboWOoRoUbpYQSRL0CbyecQ+5z8PsJPn3wywLetonRN
jmT3jdh03m/yqtxyibad3H+4Unn5lb5v9gYDVu7m40u77dSZ2159Jq3tqgZ0sHdZ+I9on8c7OcDd
NWN6RwjasEjFQyhs5jwGT8463H3Pq8GSE8M+Vg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
TloOuWBbnNfShv8OyPVAlDVmCuRJY0FhORehOoth2HNrOgDaOjXPrfH+h9Fp0U8Kf7371cZpzcOJ
vfaIE59tzxx0YXpyXFC8HSpnkUVitYUcWpMlTgiQQ3H10cnnB4InYX1EanNjXWiJ6xwzvtQnePVC
u9EHUusabR+0ef3NcvFey171Q88jHZvIqn/waUj1O/1rxs2j+SNaG2ARIF4MGNElwYhHOVuRuJVw
/JnNpuaITMLi2hL6TwgOH3j4B4raunUOjGMjXm1x2xHDgRcLg+vDaQ0dkGE5qoefTlJ+lnC0yBtz
ysJQto8q7SIV0zviW6SxZJ2Y7AJCVbniBgGuj+5mDGSCGjGNX03hm7NTwUYPgpWnrDr/mBV2tU47
oY5+q02Y6mo2Fnretl2knobdnF2sHdAEsGZnyzyhZeXSsDCtGd0ygzIqs0Os9tpnV1JbSGALBp/p
JmQFRjrjqC19DxUHxpJV9ma4eSiJLDCbhY/UYYnC98MAo0K/jUEJjuRw7kJgoVxQ3uW5HggD9k9+
aldec10cRfWm/VzcAH46jnEoS/iUkI/xjD81g0a6JKchWz9i57rWLxvrPVStYdzAFaSoh9jO3S7B
kOEYvixt7Z8pnylN/9ZYmDFgzPvcfK5z9OPqRTJ1W4btqF4Ov0ATGv8YFlFAJFvD8f3A5pdVUl/M
zJo+I0ND57zg2cuooMa/O0xItBo2Bb53BmQbrdyGGys8OD/UkAmY7WhacXNfpdub9bAYsKeYbo06
Oewf9n03Lvft2wREKwhZ/Gfpqy3TXrnAS+fBFc4Yp54hyG8/QBdMYvVfl3bJjAs2XrnFdAbNx1MI
VrfWNFv3PNQWr/1ErG08MkkcwoNN+Zjis81qezkYfBQBDvCL/3YB50nA3fKLJV4wW00E7ZOE5qSZ
gdYXDlDjL6RJc9x8JvwnBSQbO+Ydo3C9QcImB+RvzJMrkNEBoDoSEHOW2N73jPDjYUbzNMGKqv4M
LfoonJ4NiVbsw3SrMRH/naC5OJR6g7Rqd6HYUD4xvbLCItV/Ul8r9MnMzhB38M5+iJMCwq/Vt1GF
xtjZl6Y7lyUPyp39ovjMKIN/Asa4hSVxLtKOom4j4coOUgBILKBFBGLeY+jdHoQXDsRM5APDur7W
SYPBNYUhQ/1XJPfsupaRwvGsy/OEAGIn/+KiwMc0dLqu0lye7Aie7wG8Ve1vXA423bmjMGftEV2K
NWsiVP9HJnBN/OggQV4zmktTrY/jiaRN6WtzMd6+5L+Je0cJODlRe3JNuba/7w12+472yuQYbcZb
6BYLzY8dSC3MItaVUiHbfCQZzh9H5QMh2JadsaMI4OAAVCniRusR8XPdONHXEFMwlBdR+6PxDNrp
O9LBjx4MWfi+V5kiZzfkArO46rU4eZNym5ysLeOcLPRRvu4UoutlNVRH9lQXXFjvtstzz83KGjzJ
18iIwZyPJvOZn4QOWX/qMQDeCJp8Uq0dN2KRjt1ctwcDA/1aWSPnAX63b5WiILkSXSki9NGvCm/y
YsunQ8+feEED1l2uwyRLqtr0tj31SkkSqIMK9ygjCjpCY/oDphhC61A3Yy4fFPB0vGm0cfKwGGfq
sjjTCejmoMTwMCBbXAMXn3/e5f6pCo+FHnVm4tZnkDzOUKqe69xzhbRu43W54DUBE3OwMBuV9jus
ImiS1XzgUBoLRfPeUbkcDx5PWbvE6fBf6C0epOtdR/Wz/7hdQzsdfk4ZbbYavlejliyzp5sR3Hyh
M3ZJUPHSQ+r6Zqb/W15r2Bw1fvSWGq2vLuQJVMwM7zwf7N6N2wFexVKBjmbWDRI11RT/eIUwo5uP
AM8Q106B8XJ7HShUsK231+UJ4o/qG/D3OfWz2evwsEDvNSK+hLdIGnBCl1gzVn/namzM6OamLcNU
YjqXBhixStrAEg7q60PyfxpPGXTHoUU4LJ13AJV4sJ7URYOuw1APpzYm4BEWfh47b1vLSQKymOGI
b0frj6EjaBKcIPrI9Y9h4PCN3Am4m+mps8AiN2SD64hMdkkf4cMeb5Unk6fQuO+gNYP1/P9fm0i3
929WEWjpSebQEMX1TOl5+Wp0Hp8gc0LuXV6U7B1mEpse9ZOrNpX7Wmkv+nQZggc8wWavYwihaH2x
PSjY8khP564WQ2tHAMUfu/GWs+X7SVUy3Lz46ILrJOzL7u2CNu5hwHle95S4ul20hX6qrR4iY5wZ
1/x6fqI/zGcKyDgaDGf9vtmDHb7Bxl22biU00L5/YLlTlUqN5btZixcdeLFlJILlggSeajiYQRVf
QU/AcX29GDRDGrqLo13a1uZv5DSTEzL/XR+2d9U5YWvEEINVqVW39xZNQztqBwNApEM/iOo9n+/q
KtXyMIzGoUde0QrS0qn7O7GxZAcNR/HlBTp8+mjinD6IiAjOLP4VMcOzQRxQYjCZVym3IECg3+6A
0dkJH+kF7tNwOIL+sYmkmJa7O/YaCjbHBg1bTkIl6HXxJDG4Jlb642mkqdNFrf2B5hgrxOoFEE53
wRPVtyu+81W/Lx+d4ACFRDAaIa2WqPGd41HJVIGMSxxK23nOO09CUsAEMkX5Oms63BzLkVD1vwTS
WvSMYVzF0HcogwGdGT98uIca9qhojccBu+ueT/FtF5cUjv2Gd2/fVVwIkYKD24FcZoO5GFSjX/0g
UBUiB5o5y4dzRcvAiodl2F492efH7lZcsSOfv/+ikZY/dw6aVqaBUBJnXqMZ3t5hQeWkDhz+J3nW
J3YHUgsjHm4U+ILH+aji6a5ta6+3fBLChu86/+Vx2KvvuFLUB2+g86HZ8uOsxdm8zbaNpQ0F6sBN
phGcAFxUCpyJ1tNSxYJBmACJPTirJyIxBrozGapAFfQb86YYN1SfQ6d9wp8Z52rqOecsTUnbSJTP
g908H0ACVKhyAmKjik0mRdHY2KbHEp8w5761bDDuc0ym3ImLCZ79wnGYNgyvnrAogKNNZTFXUN1e
ze2H60AFVWY5rNxsBaNyqkw/yT9s/iyDUkgNLxO1wwJU4sFHXqmJlKPrdsUvk3GHfg+5COxRqP+j
fWosM67RgPUagnGauuvPvvEtopLYwoND6rViaSjUoBtDOUgVMLAXrvFwglByKFHDPYTbVGu+EQZO
3znGVe1rOs7JK7GQLV7R3H3HL2n79N+VOATzm/338atnVW8QzvZYI3J1CciyZ5aqakEn8hW86urR
MGd5+qbTis+pd+xCQDe/9jGAcq7ltS5cbx/RNfEW8Lq1q+/WNKRlBTzYmg7nNQBI9VsFN+CtAbXt
8T8KxZU5bJT/TWWAOzZnBIRr2ms0uC/Xu8O5YABJTq1MlscMh08Sp3yNPNhDceqYisDkMkysgXZk
zCey/IJKULg5TWOP7AxYK6AVVTKJULCyvwD2a1xDLQPDGrK26jAt6wiEf0LNnv1o6VCbwDxIvoL1
lskIdSTxUb4nISg/VdrO3oRsps7Gw1HYK+wFlecsvUJYOeR3zE29HVTPK4MPRAt8RO9z0WFLUf0q
9NwCoHvbuLaCq4tCNQe507J0d4i7xeT55jMDe3PQcRkCo2yEVz9+MVaDt8gYHo1ba8K2U06TOSuz
aFF8IlBx0RAMp1VW2l3LzteID1/TtfUpUfgb1tg8UI+jnhkcHFLVogB7VfYRc2px9bHBhlI2wkPM
glVTJ8RZ6yxb+hLUox7c1QdVVH5pC8qAjLlKPPZA2mqY7l/rWMx+7pYxMdkVkJzc6W7dSG8M5tcG
yTEeY7OSOP2JZ/PEnDZoPqD3FLdLEK6/Uknj1TgaCC8Ib0WAjmTG0ENkCgOAcqgm+SAEwBei0/A6
zGfCPUOQOfVL1ERF6+6BvX0IQ84jfcWGxmnEVXkxqUbd4oVW+rosTwf3gTvwimpU+vKpl1ikvRXU
jEeiyOOjtCJovNfMZP3jdMYF+fihgOWw067s4dZJfygMa5hlm+eenHB6dhtFwUNJofj15htmvt4z
MMnGiQnmi1bBLgxzt8qL7rX6wujTQbQeL6kZkln8wj0VoQqN+80ugVhSYJ8l8u80pljJOorZyCOZ
aCk37a0TbFNHkcw7UrSZEA3GiIij5Pnw7q+pcsKNpX6GrYDOY/9A9OyTaIjYsOYOIJ+U300tsdic
mrmXMYpnSzWNsGQo5jF+zaq09lp6e5WflSgwJxS+3SjszlDgzuU4Q+OErbXrnxzNfxXFNR8NzhA7
TIPp1HzHrl0RSAIyuEoq6UdsFzj2m0pmWdPKJ2VzSkvijA/o3oPi5AwM/UHzJyPVMM3XuV0xfeGv
2fKbnDWDstLOGD5JjoEenIgrnPomy6yUcbFrZCbvoCvW36oRcXnywjpdO3U8RnclN1WS0JdC4BBS
dUAia3s7bjbXbq5ewNzhgJb5vEQnpqlYN6AaTzNlvhkRfHfNxcoubYHlXJfJrh0br9GFUHuYfGDF
mZc2Gipeuzv2cfAuIgz0tL/SlGysaY9mJ8xUHhtRdrsI6TSia+0Y2i1Zng0rFU/9tyeqDhpA0VHd
xHvTyIsEfF65EO12dJkHqq/2przUZbY5cchlYew78zL+sk4ef0wIygCU60R1SLu86fwnYzpyAnjf
hLEqRQ0bcwGPnDQBEm5y4Cw3G6LXvKPoSe3Bt7OYg0BeTZOIH11KrI8lqMXM+JayiIrDmnP8jjf/
01PRpHOab9Vvx0x3NTZ4XIYhi9SMdEjw49CsLyi/gB5k3P99uIjwThRQ8R1KEghN1ZJ443aQQCsf
fZmNLKVPqICEAe5oAGQWR1zBRH3iHpiaaNmKvJPXfGXa3u3WjL7sw9w6XvVilbHdTYr4aQ4KDMHW
Ik5gNBzG/pjTZVGkfzD4wQ4keRMc+mpB1qcwn/JfczRD8SD3/+qiVjSiEXQln1cRDWf1VTPy6+Ia
vBf+x3lGq6HDAxP+AfKK9N1rqSk9f2HWBkqii5A2OGWpV+yzOKdChQyZH9fKw0AS863Uv3yDbHGc
qNeea+09dZUksxTIr75tBgTnuWXeUXkvM0SS/yOurk7qMadj7BTTyjCXON6BQgsDCse3S59I6i9c
J4kql2L2f0Ipjx2VCq9xl51+JQgCCHn5ZMo8hRk5fgq+qVCUKLbz5Iun/76bpPb9QIJ0BneqzNh4
7uajeEpUF8M7FF5dkPHrbzm/s1h9NWq6hO4XrBqGgW3Du33ddfXCI+vnUbFxVelUVFXkovDufq2v
bLU/PxBrPG/4I5HYsBM9iyCytYQkcoh+vXhBAAGJJ9FibYCivKQj4X9skfkaZyx8qyerj+243ptV
BkIWG9HgkeUOzKgYAY72t0qKlvVvZdVd6iPLwnjF6lpkv1bDS0Z8z3VeYePwms0OePSRee5m465I
y0ZFTf+PFzrjty7Y6ho8x5I31M3v5yM8tw2uM2z53GHwCDBFlwTJtXvBf6dWxglg/cPa7iYdCnzM
GtwJegrD2+NLb02Bs60jlggnAM9WpKETS9b/ierC0hOLzPsb31xjqT8OEfjLxeLUpxKJVkfuOfL7
K3Tc+NhbiOlUSdrom911tutfSlVDNOkoF53TBXdrZz9rTcpPqOL8WunxcaeOnoPGgdCJXi+BcR2V
NL0GWM519H4E/sOBb98poequClT6DkmdpRuGp9Nt29xZPuUGhM8ZbHtHR0hwX/j4rwM2xEHxhGKK
rLG1nTmAq/sc9MmI1b4EKRPhL/ju0aZ+iFuFivfi8/8XgMzFBd83OBBleJjnDcYzkE1qh1EyCQuL
dj8chKQ/0U3pbTYJjIVPQKxgFPVE02mcI15PG0yFScEAeCH+GNJUqgK3c7KybgdUzSLYB4A3Bnfm
SaM5giGlbstCcb3iedNiwT2i7Uf+P/byep2YRcYFOAZtllv2+ESm8jBs7aM/qQfkjI0RxuepQnjl
lTB4nOLx0TG2WSFm+mixZWbqtdK8QqkYB7PJYCkYt7NDa//edDl4G+ICNhJomHjwtYz0gCQTmKDz
vhJ6bb4HKQyFwoNy2olyCsHz4rlv5xxZqiIXHbo9bfwDFhfkbmtatxsEkESDliS2T+J8Bt5kHZaZ
eTaM7RhMcLjvavTpGz2KeZ72kYIz8VYYHof898JJsk6WDdU9q8Qoz5nwN/gp7mnSqAr8cGbx34G5
U/PN1E/ROdo/Imc5IXD3fNzguUWulJeguavB3jT2PKP8cGou4F2CBnj0N2jGYlNrQbgA5UQOpwSm
bUHbqZRDS4MT6B5G6SDY3yDpo4ROkpfgkZ+Ph0ekOCIwbcFcqc3I2v8wwBZm4fyhdulmaTRuOASw
z9UD2IVu4FXL7lEk+2eVSl90omGN98WkgCGdDrLLpqNhizd1hkaffMn8gF/jcDvtnD2TAU9zaRFV
5jAyDEPZil1SBxDUEWzdVpFv5m6LS4t3f6hWlm2QHTRZBeqkR+CiDYOUJHCSILVGQ7TApdEDI5r/
E7Hpgs7cquGqVI+UiA2VdK6SimbT1SQOSGkSLxy2y2dlC+8SNMX57ZaZHfZe2BTMwiK7rsjleefi
DuWtO+Qimf97Cqcrxg3bXX5ItjSZBwg90S1ZUtZq/8qYEhMv2w8ChDm7DvqYllMGHqmA7a8EWlMq
NswuckDLg1ULY+jwnb1uBHuQC2HK1S7BhK9aC6zeVOoFSxrms/F0dFo3g5HpyhZLXaCpAT05iPFu
VvsIk+baKu7R838COOqxTy9t2OFT8NQz12UEDMTEelybwzZaHqdYN3X3W2Frrgg7xUumaFNqre6g
NRCH45H/q/rDzCX1/89VX0silB/UByL7ovdPlFHLxYj2xT16VuxIY1DS6nwAhilDY00AwMbUdc6m
b/BS0GuiE2C3H3t+ROJtxNsfydiulYM5p7EaazT5NBU3+IDfAV9addCY9oFOGB+1qEe9C9/ZAn/h
+oegp5TyqtazUQOYzEGjPxOBuW0xU9OHUj8e/4nerJ5nVoEdUnPtUobB2VvvJCh8vKCLZSRTQn0P
DMjURrfJXxJd5Cw1qhzAMck4JJI1G+zw19CUcByZTtdZyudQ3/ivaWO6ZLZNy8XOCTFjMoKEgP1/
wYYlcHod2bVvh1ttPpUiZbDPELWfI9HhspECvBDKwQyzSCsKzjpwUCAlvXzAdTIeItb6SaStNr1K
SWGYwtTzxhUkfWqIf69BZMyiG6Xw0WBPv5xwNqj6mdcG21DdcFVcFkHVx2EuxPhpCdCVzzrJ6DeL
5NiOrcKh9gbOSnDbEFUZ6Ke8ZBJGsATIsiefw/CE2WCqsf3oMW6tzNxdXhyjEWLLrHTxw1n+4sWs
urQYCkl/vv5v+TubsdrQYcnx2Vf8rvwZyY6lJXjycq3BXcu2pLS54pXaCpe3/cPsMN/bu7JLbZn4
ENDdbkHH5fabYJQNZxQqrAM3UrQzR5a/UVD84bNfC91Vgm9OFYYJKo+3lbPnVbVBKOyA8ZjeWiVf
acm45NdIUU74qUt1ggXfkuJJIIZDKw3KXJBnWEhsLymub4ahM/a75pPdp/ByiBAth0d1KHBl8E/1
JyKlD4MOqlzcM9IjpNSSsNPxkB9s4lcnW6VLsWoACwHXMSxxVV1kqChNat7FxR4+7lhJlJnrEo1e
vt2rDfYK9H4Qz3C+PV6CIe/Ww4bW62uBHzr2++6GDUamvpVFZLpW/8sONr4r9hvIrzl92ScVEbK3
KQQWMjL/Jt2V0s1/UKgRo22CtRqq0SBHRgNdm6gcF46sgTIfus9mv+im8/0bs6aj+8DJDYf4fEWe
glffsjfPoBDbGOiPagYXBIVvktbejvwgJ3W5RLQ43tEW4AyyD2kh6jrMAUpFzhQ1iuQCMwJUNX/K
EVAj1fTmNeXJnPfIYSvFJBEuh/sb2YTxtBv8QBzTLm0E/rUXKYcNFp7YYh+Hmh66sWjoBORxfG83
hJ0/yg8hhqcYILXBrmxYS6YMMOfiC7WyP1hSfzFoXPStzNaRX0diCvIZa1hDZtqRMD3udjdnLWg1
nJE6RhKgUiq/jdGerXwUBC1pATIRCdPBlgyDcx9R18cDTrZMATueE+L9waO8/6bNQslLXL88lggY
Ll/2ndHtvKeCPvTeNiumwdwv7i2F4Uxn6qZXxtQKfIRPJmKvEux2a89d/bvDTIRAhx1gt3kMIRKd
uNmy0XYSkjqwQzfQMidNv72dHVeojBAEVX2ExbNwyaN1yCnlba7nQT1w16Z0DyUR5UFTEn9ZQvfT
cmssw4LcRMkAI4C3whNLKXRiMdio+JHl+tmQXSiLgQNpLwLXfZU4qLOGftRjmLJFm/odIMXEaMgL
fbIfyavmnS1uYPwVvh5dlwzg4QGP8I6A79bBnXo5F+eVDTunWH2EZrHXNwRA+7OgQQBO8Y5O4upZ
I7KH4+gWolp2u7XOIf4NInQejf/zFlpuPcf2kNQGsvPkpAqTg1CU0sFeHIh6COflIJPAGrXea6d2
2VlwPCZZqbGxL1H5OCNrwHNHcPxcI6QnWcSrnzRcyOkWJp/imtpzSYFIL63aDHC3bZD1VYhbeRrd
vqnPMl5DRedFnoipZbscNDxTfgsx9zXI8U5jzKNENeEoZcyWCZjdkzm4IBlymZOcP9jB/2iAfHZk
1u/3Cyk6gww3t2IyPl+ICN7n8mGcJFpWS0y3QmKdOqAV6Hs4XtdfAROObcYraCbdQgahkyzLKhsN
sEhOBB7eT2BdHvLtffj5i+PgO0Cv92jdxWS888GZdgCVgZM+llupmCbDRFsgW10cgngOTrO+elNC
CG2dwYW5jTn6iwFZ0auoRtZwGfnd5vwWIDH8sssd9sTU+YINuIOSoL/pO7xR2OyPsFZEzeSez8XJ
xR5Q8pPfcQ1q2jKOmrYsg7e6fpK1nFK/ZylI1UEFZffddN0NTFIdOscEM/oN7dc5MOkhw4jKajZz
AcJXtgeETiY2+E2hH+Sj4FAuUGkRIITJ9Om6wgoIRVU6j4BwTUSJoi8RkXaRgMUHG8J+CJi7T/ld
F7ptJuPd7QZBVGkUP6TDNp997/00qTrFIxPT7FUvDd4i978Xrdc0uQ78CG0HYYXOOfcPgjSL2Oh9
oE2ixzJMTZIgun4sPxvk30Xn/ymlLpXhGkX6/XtvdpET4F9xquMEW3TgCYdKCcwdYK1acs6erXvz
aZuNd0njs9LPP2Sl3GFW5gYoCfnepm2KZkHliUvYcyRYrMMmknL70VgwPnHIyrMMyhEJleWmittf
jmrw3ho4ol7eYeq5ZsOK5aW94bE/g5EkTQL69RSok1ZGfjWLpZSdEkMosKcvHzGX8wWnHsFrIpZj
LpcofrOJW/EXwYqeKLkY7Bva/1gzzeH7seEoS654QBM+hv1KDeG7Zr2gv1+viqUp5cfOUvNxogFS
0uxo/7xzBVuBoSlT1wBKOhziS/IgvFIN4JlM2LMOT+unKyiPWlkC4+q2mLG1MD4TJ62fT9z4/XkR
4h3iAhrizBOZ43gvOq2Qfbg2qQZa6m9uCAbeuLA7u8/nrbloUVqA0sFF3WyVtHD+PU2SIEzTq6kv
WS5zjmLniGPxv3p/6OTT8LLlyQbQ8rZw+NK5MObxTj1qtbtm2IL3PtX8G9/e8+VeI7zuOh4CqLs3
ZGMq9dnVjCqlhSerRS0xTtUl43nMurGr4QM8PMWWY18lgoasdjTHDFRh3L7YwmwKurwLr0K1r7VB
2LZsnb/uij9EKX1FQEDJ9C5Yl51rV6Q52vgkku54APcPAowUnCOFmsXAnt/tzlK42bLYrDAOteWB
WFVrWuR+k9RQdSfX9vcL3a9c/fK6K+OtxejwUfOfAwXVR56fSkCf2+LglPjkRQEt9ukfYOxJdjMY
PmNZGtPU7whPLeC3tAkpfc+LN8gxcS9omjGv7BUT+ldkrH9FwxNWyvaf3WWsXa1piHAiLS8gQLYA
vJChhTjwAW1l2b0jcZUVj5jU/DJlBzM+mit0jB5ozrcWajaUeQro3+eLrGkV4G5YvFmqM6hIfc6R
2hR1n+wgage38siOYAOe4MmoOHBYWc6RT92Lv/gQPvz9lOi5QhA6x/weXbOon2vc2u2YBbZcQAzk
+LEVnZ2Z4srLzWfIcJiU0kA8mFsvxoi6JF7eIf/86h5iPtPNpU274G1WDpT4/aZppnsS6JNFfNwQ
kiqMsU3xzSWcAZP/m2TsJ1HhpoEuIVvoAevTiuR/y1ZsqHamfvNtG/fYbtJmbLKGm/6jBRFbLp8Q
BAUeVnliWpybcGY6sq6l5vYbsngoItpxWie1GYVxzyJXZN2VNcVWeYjMFg1M/H6b6GJ7AHdvon6n
CB3RCFf1EvQdcVm5i3yTUY0aFqDPbQ+a/Xm3s67Okpf6izrwmxWPeogwaT9xl3adeRRkigAPrDEA
BCfZcQ5W93rQ3ItBQyaUA59nuvd3yf2EBHYyy8K9J3Sgm8RXJidsfUWXkFj4IwHcNKAOYodKrPl2
lUCYXqZyRMasj6j226K+mceoeFLTp2ph5XlxGBamM6V7g1Cq3ljHwdvyMgdqlVbG5WxR0dpj63N2
zuRfsJeolado4q4ndvXj+O1isaH+nxUGar7/KNme6gGYsYa+V4wzV/t02UVag3/sAFr/ZQslmHza
rrS2Cl48ss4/mUHcXwREjP1ZVT1xcoRRjNcW8eqO+QqQOImPcHgapKCMaYK+J/Xe2lU0jQOYRMzt
TlsXS/Wdy0uMGw1Z/R2As6R1QTnq44B6IFoaZRfZayjyTPGovGyWm6314PJ1tCGaZIvD+KMy00bj
s/mV5wDQC5ESVYG0SePbCaP4zMtenVMMzejyAvqtdVDAeHUKzqOTnkWDDZeAHXlWzDZkpPLD2fkK
ev5uf9PwM5rEYvfx+v/6ejUPaczdorOj3Z5WBxLq2fbI+Kc5TLePW9nNDUNooHo5O7wAfkkuXbFx
tLh5PCxV/FL2jXA25zUb3x0V0eVdHLlAudzXK7XxjZQPpp5sEhY3/4OhwC4ASWFmgEHI1LzK79EJ
ZkPHSnCNmSNWSZLWc2HhpIpeC4H7f3LjzymEtF+aalBvh34pG/zfXYF/qjiAUA0qxuAZVcn8p6LR
ToL83ND3jvBp8GkJJkeXePfkQkWpsby9rxRiZJHS8zWU6/qMIhJb3jaPVV9E6VF7cEiRSTHsMxGb
Q5n5lpT0GzwMn5bFHofU8x8eIoBMKwCJqUtK15rD0Q4wzxliuexFwSRCT6pcp5B0sFWJB/Ypktmo
lVXSHb8pWX/xLWZSK2S/fu7PygJW6wyXVDLt8EAou+UPnYmU4HeAjJiHgzQU+1bEcrh/KN3/UzTE
gGFB8IWMcYf0gIKUPVoBIngr19Gic6ap09PpuDhZJoVtOV4php1UMH6hgYgDqLzCy+ZjwB2MTUDO
/i3lwFDYwY7YgsTVp0PwaOC41nAPRqK3jToZ/mHkxpzeSVggOupmecjoS3bU7s3ZJW1NyPnLa2OO
qvGHZmTjbEnIfB+QzgUoo3c3BGZ/sEHo62trBbOugPX7isyAiY58z/DxaNao2W0bXNE0VB/HlkRp
Uck9D2fPLA+tynfDIE+JNnK2aJ9x5Ren41hO5DtcqwTEbcn9LZK4lXE+QfoUjRQ/AFxXdUQL+jow
m/8NdGPt/awjn0NAsXkWt4TbiPAAHd8WIR6p8a33RRBPDP2G76+H1QCNotBXO/sZcGaFCj7l6hUd
/Cady6tHq7g6NlikvmivQO0kupwD/NYP1qUt6oAxRra73OuNYByvVvzZJxp7NojiNlohkrxeqS7U
lEU7H6RP3zbKnjg4dGns8AbswlCflH/PZaQwFFVGBDl5qjWjg6ZTspQXPbqfX+ePMfmk1Pf5FYGe
iCouaevmEDAoNGdvEKYS9KzPciLsxXwtc2ExSTlnLJ1SIrLOZTdU5Q1bvIb/E76MFQcTSw6zOx5c
DOiIj94/ctRC+cNh6jT5OqRK1S92oydiyyKIq4BaXAdjzyOMja6RFswN8jRqWE18zKEdNjFULBN1
7IXesjCtS1q7JcbW8j2aZwIz+AuVAbMiA4tz4dCQHF0+VldC1miaCS2Aw1Y3P0PCiDACHJ9BUz0q
xbpv/td161BqEwYyF6PgJLS87gVETN1QBOBtphyjvYMVVM9ipBxOEjvfD6BaHSvW2olGmeyvm4he
L3n9ShDTHQOLpq0VGE9DDhPTM3We1ZCGAvcLg2iNamMIrATkrF7giSd5SUjPDMQGlgsDdPnoVZmw
pV5evdmgwkN7/AA9J2gYR03ux76uoBXx0mt58O+PkgGiWZ2VRsjLCjXUx63T/9VccUKvJVeYA4E1
JIw+1DLRbXF1OAUqwcvH14FlPr0k9G2kQxLO9SAxcvp0gxppj/BdJ0/yi9OX6w35r5DZtmfAO9PR
e8T1minfxaThv9BqFwJuJUiDXpynjHYiOtFjUhxZSVWk51mHGaWc1tPhqEb6zQnusQU3G1LMnNOG
fxKfgqVi+4p0CdG40MbxPORWehyBFeeOiZNuS+WXVySkue3cosqkcdPttXjTwg9Gz8r5FaZZLSmy
TMCbFuIJqqVtqTlrZ5zTL4RHUGP1kzKtWdlw3wlZTQKEJdljPyCtxJqFX9rcFE4s2WGBHTdu7Moo
JNhVITE3oFObRfo6FKyH+YkMyQ7AqzFotNK4jPnC4LmmKWduGLjSeuVss/6cfitxoVAVAS1rHqxo
Hz/6wmP+2zmMfzYjVVPksr3zE0nhJvPMXnH7B/VaFo7sNmxVP2bpZ7dQJsbPy/AlFimfjGWOj3BR
gF2ohthwkTEHg45cdj0r56IRIUzAKTUSnSzkRn6u0ygStW3Z1Be+FJzjobrnvOTuZwH4YRDJmMlP
mvsLqQtVi7+72qNrJf/REl7xk7LfSs9CE1EPEArqVjtiR5UNukMSHEVMhwbD6z7uCsycV05wKZ0U
cnq20pzXpeUYcMqL2XcBmDiUGUf2W+22VTvw2jtl1GxDO2W/sTuM34Dh+DcJyp+0UjEgYHaEeUBr
dBxFRwkkgME+hJvYEsa9QaZWkHGUc4Qa1/2NlIHVmT5m/B8SGF4s9cSeH3SLmrMglXlQ0qEYjPvv
+U5aXOynTLCxd9Rg4eNK4hmjVyPlEFbvdtJNNeE0W/UIl3LLoM/4/g8nWb0JWRQEC2DnF17ItP3b
o0zI8l6IFvdIqujZqo77G2PQ81kN2SKZmlPtHWrFsdWuCLIBn7wRo09ba1EI1Zoh5SmTUTfqPGuG
96Jt6aWUwqOm4zfTbUKmNuwirW497AG3/2RFcOyGzYKN47QNPwt72kPJRP1hi7q5oz+PgnfLLSnS
xUqw7pNszVEIubeHH1v10OXyCygUaWYyJtX5xBb8+PfKNlsA4aiBikUNeZl8ej7OwvfnobMkn3Li
VKljNDd+59bf/1tufIiVwfUMgLt57CGrE97gmPc/yCrzHIXGItjfC77hR2fulq8/YkNVa9Iv0uYA
G3YgRvO7BOlC4NDOQly4JHZdVFgWZZB0BfJ+1pby72fm6hUjbHzAzbOQNl862rYh8nWAG2rpL4u4
nW6b2aIQrSJ7L5RIXG90VBTXgS/xJnoXGeEFgZ/aZW/k+waBXNrounq4eTvExT8crQ2+0wrTOjU1
G/1lPL7v3AYFNdx/aHDeGja0U5LghH4l9TG8A1aWL2U6irxwLGIqiE2Dp/vW7KOhRfvp2oUrPHvZ
bacGWxQTGu5pAw1wAQBuYNplR75IUWKQBn5RO6fJJsaSPtqsbTONVCapAltlso36zMoEIXvgdjIp
0/+WL6NL7auZURs7TrGLVRDfwjgHc29ocymVlfrI9sGEOoXcWMjQhjoC9vuvP7encl6nbORvCNU+
mcOnLq3YcAZoc1ajvvBQ8ZkLmjnEY6zwdauTWfEZicWsJWNB109OMgHTyMXoUBDk+jPFLY/s0eZ/
l0Rs2FRPPZnGJRfhr+09trMaR8CtCCx7AXN7lJeo/eYk72Py/Xtstt9z5sI/jFdmNgWpClpgpTkD
HQb6t/BjhkqRw7KCXDH5g8niPGMbPCEcXp6NM5erbceLFiPTtywktUnb5wbUBZiXAlZXRokIiiXr
So4jvAMcWPGYGOwmS2pnHs2o0HjgCkAQvSsTQR5XWrDDgie0Wet+DjBVUM38PT2S0WPBgDFdb9vo
IakoTrtElf8B1/Sdo8DyOz1l8V9xOtbLwTORPJFZNmWRzT3YHta190CLOFFnvZBSURpqrnZ8kQ1U
hY9jQNeo4/cuks80yOMucsnfMR+L8pOKAy2SEND+4VychPonc2LrSNnGk1tsXUjRwAUVxGR0QyQS
0H2GKfRjGkYrrwFrCqJPUHU82OL3CgC4I3BoAgl6LQrBrP1pOFTWMHax3xQzmjaW8a//LF4tTU1G
JRQVyxXW8tAfF0m+lDVw0phtqce4QaTnFIj5slhmlkjhDbyFKlaHSqd1URxXH5ksTGOlEH6GgcEE
NIfM4MP208lW04UjiYD1+YKWpFQhga41BRgK7ztfksHieuoBtXV+J4xLaqylf5L13R4r6b0iK3Q1
l97jA1V0BKR8E+giBk0834tDb1EObGs3sybcen8vHf5GWV1IRjlE5PFLxNemGMm+6VbQuK7frj4V
sn8UVrwZJZ8N346kX/WsERwLvZ72GcFVKkamENZwxXOLtvoDf+yC/bfxWly8LJHnw9/tD2eXJ/ZL
qh1I7OZEXLwbrDqRCvmlP6ybeeb5P/7bC42bGMMc3S5PF46cZSBAE9OGOKIbQfCvMnosxd4C1G6b
pZ9c/0RPXr1dCg341YAZNFDx3bbEow1okmBcukCb+s3YCY6J/4kOeRiL5YFnNC2jqxYdpsm7WeqP
8hAHU+8XyITMd0JXpWhS3mQAuXGTGGQ47rtQCet5FaPdV90BzoX/39MiLeXjRv9xY7YBI4P8T8Ap
hL/t1gGGQ5bvlG0xkD72rwOZsebHsEB5hIYnXHi4F3q+DTIRUVnKJltOda2yN99SJxICRql97ejR
O8U9BNM=
`pragma protect end_protected
