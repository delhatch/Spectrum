-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UNtpCBjLsqb2qPQ2bGlmrbh2WJM8YrNxEkg13hwant8LcwR92X531lM1iPucwnzuPTT4v6eXmfQV
bA6P3Vq25D9GFIXs/TLxeq5iIBhG+KAiX9F5ERu0pJyQy8ej4HOcqAQcA/yQx1zTVsohvPGcvf6/
dKjdNUvt7iFxsj4tNTjT/1klNo9lE3/tXH503PVYo2iX8weh097Iz97AohXIALyIplN7B6XWbpQA
FQ+Ba0Ni9I2T8nnCuonQKAjugi+2Z/+GaF/tCoX2e9MNapswgsnfpRs/oFCTnLFGNSqjrmkQgD3i
6o4d7XIEi/9T7uQhiGf0IIMqTryUaL5kAbg+Ng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
x3YNGiIokpVgJh2godbUySXzncYJk+bk5vNbi+9e/vzjFy2p/Lv4nAZaIS3+J8tDwtpjyMTbiPJ0
B02blvoFb2FBpS35V8QQ1yQrdD0KABSCOeDn2rFDqclG75xf1bVeflNR23dJKXn1N96Bo9eaXfUa
ks/OMvskEAnHrJk7S+g/ZlxACZztZ3KeA41tuKNh837ddQEBO2Pzkkw/GgCojMWnLdeYiNwQ5WXQ
OYTN0O7VDwAm/T5aVbOSPAR4R/299s/mPy+4g08FyobVv7b4V2GKrhFEBg84ABhEs20bw0cDfM6b
cCh/c9HTRVKP83r1WnoD9V3At7YfbbjY0075NJuIBPFRXkkD5A/lvFgJjy3KdbajgkaVrkeq79fD
DQ1j9BcfaFSTMlv0X+xTirGq03Pkoufanwgudn0Z8Nl9A7mMhkhYv1mkHF5TRIhVmaw+XUJfAvQg
1pj+lYXOnR3ScBEJd6VpXONK9dZMl5Jch7lsKwIFVXQPiOZ09xm3a4RWdJGSnOoD6gCvRkYh+sZd
+3I6yB+9p7+WWOTJlV8Y9Htfb/ixx8ttA+7l+2CeJRuGMS08M09goJlLICzm5CLIXpR+mSun6rCu
RTdHcTJbCwj36qhMzkNjf9PD2Fk2q/XQNboD4amlYuAORR+jlp0UCE2YI1mgPQv0a9gDNr9ic0Jn
6dTstsOOlkJNktCUNJryooUM6IPkbmIA9mFAtJE+CqGaJTENThGl+Q2yQuf5H592zxdUuKh1Mumn
rkA3umjni0JTCLCXSxZ589RpEKwbngq7K0jjuwmobjOfKKF2wbDAIkx6RvFNQmgzZZuu4RTnlV5M
KVErAZ9kntq53uGJTQiklXlzDKoQmt+2UesqEl6fefv7XhXHvB+mn7HC4rxkYrJd7E2OGXffrQNy
l5T4GwRPj2Ss4r0k+ddp5CPyWDIJCJhywN8vN29SLV0CwawV5tBnnQNQtAKeLOvRkc4gKp2hPSZl
LO5dn1aEGY4C9i+atEah/o2q2S/+/kYJH0LF6giq0PFEnxUlcEM1rQuH5j2YH3lb8EyFsrj6YHS6
oOYGANECCVmzZLvydFQvBQ2sb5Pfp9VsmgK8FxTCZyr9dquwwmrWl3dFCYmWjS0XH/WDHuLNYU7v
g9MmygBWrYHrIC5C5sFlYKCNZgfyk+4gj5t7qq6yGNEHQ8CoP8j2qCyr6rIn8hcad8Xob4wkvNmh
wxPTKTXEhtvIXAbTXTbtIEchX3arx1OoAsj3eceIFoRFG136Gzv5odw08ukwttO3Ec653FTxTNip
k5ACmZw0BsxJrrGINRUEAWjrYNl/cUSgVv6Co3EUggs2BanQCj40zxiKnJipbBuyFcQaCxUSEh4O
+nZ68e6Tmwg8G+GVEhQcyVY/uUHQry0Sv8ZkmDi1n+bNQk0GWba8TIMz+7nVwCpyFPFValVvTS1F
pf7oO72iP9mPrjQfDIaqPr8mLpvAonMoY7sLHv76AwFl3I1BnDNv448esylggmkKdO0/C4u1n18I
EpTi631x9CWVpmHv1+c8HC/uehM2s9jo9DKQDrgF4whNpYKnQUF7Cq/cSaA/xi0v+xDaIF8bVMKr
m1kVx4ySUGtRvigyrpwAyImO7+bXv2AZ7y8ME6ZisgBTSfWZx156jgX/EsZKqdoWT8kkIvwnuY2L
TF1f2B/x5wk6p+33sHYhE6Kj86pXyqbNeFBOHkrc3L+y1PJs/cImGjfuCJ6ThT+nP27nsRN8buSJ
y99s73Y3pxrOOVsmQE8OoHBJuv4WfUfY8WBSGvLe/ZZN9DE2U8O3sv5AlOG2Q/wJEY+f/67oPVU1
ZQ6e+PAd9wVwlS/EBTfnBkXpz5AxdXOInMq/xqQqlBphfXGEWhe2/2lOU07MSgevMa5sa/Ssv9zZ
yftZFj8VJDJ4/Fph9kkTepaM3FVBxqpLbI8qjEa/dA/PbSfrMshumSwDZMKisB4ijK9yTDrg39Ba
Y6SUZQXvJFi9XBZ7eMUUkQiQBrtIZKzC7Mua+DgtH88e/VoMjt0l9Zq2xqvGyry2P6kEXU+hWXl9
x5EspK/44hpBZxN0ejndlSAfGZ1JIp5wHNOsiMutvL/lykev4Z7hi08hfZzWfanjmb0ev1eOhVkO
ww3tg7+2qzCBIRKF/jPTyhJEq/hSRS3CVjkRm1Yw6ObS3ch8LXHTvJus1kKWvVP05y7yxqr9w22V
NvhmfqQO4iC3RwfFIYbTa13XZEWsC8MCnSPChggLWplAVYVVnYKODccfKZv/PW7wo4TcAXPn9cB8
qOOj/JAvlW9thIR8CDWitwzk/xyC+3N/zxeMpCrZhfFQCgSAcayAutYnO6SmEWwV/6gKOapTlcVK
IyMtbhE4M7aa57pCmQ2P/JrwgtgKgas+KCKprgyiXkVW94hc9KRD5cetzOsKJgthbdZxIGIioXNk
J6kLPBJZU/iurAyN1iacP9JlTrrzzT2f3MRQd+VoWN2gC+ZSOjEh1CP+V53h5Kxd1RGV1l58zzt6
EbXv4H5B8taVttyHiKP1soxv15Dp+64P3O9dh1rIbrft4XRIzpfJngH4Ir1v97EAMe+NJHBBYXw2
jv0/Kqk1+ACmkw5QKUltJxymJsc7RA4y6LAjOHpBchtVWEUqm5jD3hj9W5gNTkb/iByF/F0VtEVA
PKHrlUVVyjHnAVFA+Ak9EwUEIZHLwX0bZvsLzIE1Z63o+9g4MOvP694GsfepWYGO8Gw1qELdwFQi
I6iMM9EQ00yaeoNcdZoEljgOtPG2m3MW2skCyRwn8E8lVECvM3xhbZDYwiQdgy8MC9+EEyJ8OsTv
Vsa2TeOcIYDjczQ6n/tYM3etYbQQ9ufyAzXTFP1CI64zq5w7ADk+1ZgAW20SQyHbEOu7c9LOeys6
/e6JzlieZOOcJqKJK9OT0vcnI9p3n/Y3TUeFXJEWKLtUm3ry7+xBxT2cWDwOH3BBne+WR15EZR8W
pTLK1nmr1/dOsLAhyHQ3nFewejU1Rtzh66VnQdlapjRbGRpaIYhxECXkeY14KXnzUYy0I9vydLFT
M8CIFUwemmXpDjmDjy4gTxtSL706bRQJa5sj1nO3WGTDXUbNLLTLQ34Eb+WRjsBE4pRMMwa/C06q
UFRdct4JEYeVxOQpVE+CNq7UtZMYfVlKbUMl3RN6tQVJkIhV0HKWgqZuBoQV8YQ4OjYBET/OO0Dn
SSUcxEPdnopgzLu6nwSMWlBObdVXwixSLyCFWv5v+bWow2ugT75Iq6TKGY3bCJ2/GAmEyJ69uwVt
qywpSYCamHsuVefEPO/Mh/tAyxkz7mUOM3MD4d6BAEtnjQKsJDpbMPL0R6EcHslk3HaS1CRaq85N
xTPamY+mkI8/eDEFpZw3osEen79wP3QzR7IkIPa+cYxZW0NtymaG7f8elwKKchBYmA6gokgBI9/4
V37ZLq5J+fwlsMrDntG0+D2hy70+bec8BUXEh4r0qR1CqAdDjIO+rFLJ3lpwLB0kpNHqtUpsMoJW
AmGSX7a5q492uan7EyVx6BYw6X30Ao3BIjKxc5r8t3XHkw7PJBLJCZLDCrTzW4w5D9jJOJ2XbTaT
14uiD3jbbL9AOavfHVGBPVl6tatNSQCn1R1ceOQSxnGNEvxA9AOXsYRA4rNAdLXYOcKu7oy90+2W
sEyjnBLwIRxNJ13yN1gUv+gi/yPoxrIt6xq4mca8a5FiKOhWQ9bgV6Ha0YFxSlLs3JsZ0Gf8r9cY
G/hkjU1R7U3XxU6moyNVkRsFdRc6CyFrD/7+dUuh6b0cc442r9hMcZOXqyQQr6YVT1dO5dBsIDzF
YvasTQ4J6CXT1uKxVp5X7GlacRU7aIdNf90YGSsCf49pq1HcRBpHK9DLsOL6WCWCrdTxB+h/+4qx
10HY3R/6ZMdQNeB2LiM331w/9Mv1dmgC5xiyZPVt95XTtvCw1I2QiHl4szkQjzziGydzx/krYmVo
tsru+WZL0FTx2WYHridjwxVqNJMzaQkawSwDu4+QJ84FSzcBnu+ggHBHELn3RkhwLtraAxjLejtW
ZjjodbwnthQ+o3B4YEmdAMzul3XknyqnLVatBoSpBEO6QVEotPHhuSsfBH0wdXxlUWyKAi+HyRto
L/pOO1G0+9M0sSFIMwoqIfSqB/EJFuwRfiL0p3ycYxzGOA/ulB3OsZfg7eDXri+ztz6YHYHFqG0u
y8fohkbZofaJQr7jM2S76Zp4ZMsbHJHlOCch4b42dZvWW6yxZ3DM6Hoc88UPe2R7xL03kM/5QRXq
xg2wo1vv+I7HgTJxyCDAsX1vR//OX4Hx9PHypFiOiGiZoDoDoEFbdhShzTc8ikU0ScAQiG56F0oj
MTqczn/xh4I6Y8bO5juOQRdySXynkcB6CCVNnjwSpLRSGR9jkHYUGi8gIoG5tzAXXSVgDvgYYO0c
/H20K/xLLpYnUa04SYNDDtnF3PfgRbDmyBjmXJjad7U8syt+jAbVIt/FgHZv1QbrcDLfNPGE6cyf
X6OzPbxQs1ziYaqynsldoFIUk9xgzXVILmYGcSbou7u1GUP8SRa1tZZW6zBCN3cVT0HdHB9a9d4X
mmODmNQcfh9iGvVBb/VS6DgtOnfYRNmusURSPQAgCkppSdKCfSX3qR4e+h1jMZXoWo2CGkUp9Dsa
qvu0MmTSZ+T2dV7Xk7TykBy4qR5b82lVLeATgw6tbM1kZrQ3bne59WdTNxmdlXt3Kps95BEeVIpa
SKapCvvJnZCuDwWLxz3pkAt0iei2nPgOE8zm5eF3lDpNzjcJ8wwPTxnWZi/Lly6Rv4JrKBZsUMp4
krOHpSqjkMw9hElA2zLmnYRKUAAW6/aGEz8JCgjiVV9Us4U71a5hDeJ/CPYQhosMAm3B6FIW22X+
jwxCKuloTq2mIFFlMR+BNXmKGl5FqWgYr3M4NQlSRI169KQEImgTIp6CK2RzPJhgncqk/lnFaLMx
2Lm5lbTelaMQ5zLT4oNPfQi4FPcnlnLuBLdQzvqLjo9U7T7+xiND1oAaBsqg7uXGGMsk1tKeRpiB
pX7ekBi2jzr14Fv/mC9o/X3/lQA8kHfQSt6+Uutq9kEvUoQBOMlHdJ9A8tFNUVeg3X39Qg1JikOO
1oVKpzUOrX8R21adN/ahgIYhDUAWKXN2HcxX30q0ZiARwRQw36ExB4DAX0XiRA1EFtFbQ4+s7IHj
1iRyiDxepILhK9G+e2oU617BtToJAgB+WgYm9afDgcBpbLeVBcGldMKkxUVlPgPKCJ7//qlwehZa
ZHqeuAOvskXNQWq7J1BHpqefsQOCYd73+ThA67R7Hgf1WM/lfWrkp/GZlK0FPI5iohJZs22wBlhv
ENch08MEsMOBbZhpJxzyYDNYWsMpm+3B3O0DIMBX4yIcv4SULjP8JrAC8SVyvgwOVpokV7pR/N6W
GIMgaiptFjYoA9iYxEMTZaYyusWdzBvm3qCd+9d+9gczt+/Y7zpDLtvXtflvARiJw8FerfUgbu/O
UuM2lj2n5v4Qu98S8PHjG295biGNQAgHLiHo3GPR5Gh0fDOb0qsf5HSuA0Gq734C81xmRjMmdo8b
9iUKq8uokCLQZUNCin70K93NHZh9nRPuFKPr2RK/gFsaOmcvMDsGcpOu9o+SY5c8w7mhWGAWDLQL
NAVI+n5/LtonDZrMM7SeLuNCiJUwm7/hMpD7quHiX/TwRImOCXaJ65f/6tChWqdL9rJdRbEmg/Gc
P5Hva120NZQxXzgA2XxQCV/N7FYmZGgawidTIOHsqn5SIk6QLktX90UWVbZN24hdlbnB/PbwIvqC
TToy+xGboco+pHKWto5UULaS+LQ6SoLWS1O7kBRBTA6Qp9jDVcLfCM4/CNafMWZAf+hIq4ySs9ml
3jdMUSAuJLJk4hDhQrKZayX4DRHmComzGhEMyebFc7rUNefjhuQvBVOdS7qgNgdFmqcKMRTfLXRY
H5JGuFEeU0fi1n8lOelG01lvjgopUT0NveayboMZ/t/tpT4QFQfIcaMP9Q0xCnlSkGYtG7HDOKoE
rG2Gr3e9MLiy+8m6K8sRF/VidFF8mS0C6ZKhHI2F4o0/nakh+96dkg7hLayZpnD5s5GGPZCdX8IL
/2wHQn9F86R/elE3hTWf7Dzw/NOkRnCwTfCwR8h+cKdAIT0haFb2kTeuAg3zepD3WLs+EFIJhVxn
8SnavpfAObPJLDNWJOePc6EWUE6N7hIdfsaQugmRIwW9RUgmM9I5MCJDpCEavy7B+TIsDFyIc81o
b/odtw6pVh922iUUa9oDQBWTtxe4Xp7wNdvYlJ5DcwQdBMda6z6CyiEhmp7aFL2kgsfi1pJVqYb3
tQw29FGnYZW8cRUkv32nPpGRMfPKBpa/uHsJCzWitgI76cIqUk01oqwhrHTrJpbHERwvwl6Jz+7o
uubsUOGM8kX/KBVBqJ/P4wF/gxuDDm1JBTI4Lgf8eSf3tcWGkJdzj3fbmVH1SmfDnOx++SbhhovJ
DcxahNAsQM8m144eu6Vrtk21T1vnPnslGUGppNPLci5UilmxAtGjR5uZhq/2EmPPGDEWDzVNzzbK
3R3bBrk3ql8W4Osq6gGCuUsfRR8mc1x9qwqZWCD9K4tyq9+ctOHBPAbYJw7rGIkNYl1TopNAqB3Z
lo5YXkbVN/2PVh3XAN/iaDkdfvoYMPU0SGTE+MLg0p7LA1QAaIIL66DHXBsieTCg9/K/E7+0su4p
lLDvTiNNpE8BslwpDotIRzX+MbxX2/HG5yxT20fY2cVRPq8FqMuJtrFnr74MhTuTqJ+nMaHwTdSN
FczU5uXtJcmEXWynY9R4dB5DN7zFjAFCG8kxrGdsMexvWcp3PxmOBgVwHYxWBUTV9D4fLE+ruyYm
R6mSwesu2s8C4Eu/jQJUQfCd/o1vjnXSpUtl5for1uZrCKJRI9OfFQSRbJxS90TksBrSG+M+9MqW
YqvP187G0wlBAU8DdFz1Q5nqXmk1OkIC+cuHESBTGiFQL1YISotd4fgIJIkq1qhxyv4gCVSODbMT
BwWta9Xq4rVYU1h7oOXu2ctgZpDI9U/TiNfcZnP/nxuP8ou6vAzdwqJNxMuvzVcgMATJxL5t7KHT
B2/fwL0E2dfnNAjjRw8jw9zDJVeJAzeq+d0XgKYPhqnUPsvyZf26MwSLMkMTk6l1qtv7F3ps8IKI
8fAh78Btt0yZqE9X1P6uaV4caN7rw3tlDHa631aqX9UCGN/d69Wk83aOzsLasmhfToMRQ86hChwf
W4xtKMmoVsBOhww31Qo6soTfHoh4rRHUx8yAyhReciQ5xgEx3X3mVQPZUp9k/ollnYprZD4KbQmz
mqlaoYMI0Ak01OmJt+ZZwiDrPfzslePmRdDGyYxrDi73ezNTS8TQgBqTj1eUM+L5DRQYEd4MaZ7W
87n0x8xDQbXHbZFI6Z4iznEYzZax9b4Q5V8l/DL8O6SQRW0GghaQWO8jxMAshS+DLwT3KTxUe7LW
QZyMnEC0GBHp64IWwg1GSQRXTaG+Gmg1UWHKnCNLUPY5ZaVbeb2cMSO8pQ5fHByAuX8SZusWPQa7
pwtjZEPcM27AYtOcttTKSgvPHOThFcDNnPt+iMlBP7y5q2ZBFV7/f58mUmLbE1ut3UAxuaMGK2Ad
/pQveE0YQAqAaS6HiiVqS4rekkYz9lXmO//gJCGUPQovF56zL8eLkrswdNn4iUvBVeHy9MdEsQmU
NBC5hX1UjyhR/jCcBhGuuIeKRAF2Lyd50G2DDsDdAe1wz8Rpq8xewtA8Kps4+W7Lb8NQBBiA9tJG
8QI0lGayGZGWR0SuxAEOKHfVoTQTp4aFZb2rPaZgh6jPwZ3AIKfwGHXpWzBiRN6V2MTw1yMNFMN4
qkzbLJOE/ayHC5XM59BEUnudueaiqzkOQbsEpKjpoyUcxHxuCg9nhQdvdzDzPe3wZFk886cOthbo
eoStWFDkVqABPEOZSU/q+Bhk2cIWuCpdvjZOs4Z7sx2212dxO5D7C1PJQj7CgUKwdZU86MTa/kdy
uaZC9m7GQwfHWtsamu/cvHkToin1RuIEGJiStBAkzHmxDEonR6YEwgNiPp4DqJJVqV6NTIEE8zIj
3wqdM0VzLtQ94ySEL17mErdyH6kauAkzESTvpF1jE8M7P3/6jNXW+qNoQdqDm1a2qvpEskm8A1k1
uXNVDcF7sDXioO/9u+hNJO7VBd440YYnbLPmxHUIFeBmfsNVvipdWTJgWdFPVJHBtjN50zmQSf10
TE4f59BWdzK/AhVpi2/ZTU7M9v8PulGV3CjCeBYTyr4LUfqWlcE/ER1CDUvVCBQYea1oiRokSEZX
iSFSDULYnQ9+nr2j7wjkbTVrftIMR+HoZ6d96N3Eh2HNCGIxc/t9IuxfxsCAtZeuudjkJGiyh9px
Fo3qRRW3xymJrvdKLhv9lknxZgDsT0YYmMzfdy/vI3Lowbfq+z869nyX/W3rrIVDK+kXGICzEbe9
6eoufFxJjeUn78cT+hHTKf+EUK9itR6fd/9BU40cUbm0ZrYjPfBSdp+YNO/PexB9pp9mi8G/ixa/
ljzHgX8XUag8r1ayrhZR7KMmAUFBtXgBxf/+L5cWsN/wCjkhO2bhUd8mzhIRUKTIiYin2zD32rOp
XEwVkj4sHRW/aDYT7VqQPwW4YLnERqlkYRZexZvzLtl9PDmKFsU7RPRshl2QyG5AzQYriOZUgTSY
ScNKpX5BQUfleB/u84s=
`protect end_protected
