-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
R1/p8Q70uuM8HeRWiScg7kEzyG4j1SHmQ+qKb8VDbOwkMnSBH++LlANtkaDuzBmEsBvm0btSuaDQ
LhVS+3M482lMXkIw0sFOIgtZVAQh5qQDG8ON/GUQmhY3KPP3mVNN/tCo4PsACli+vreXXl5ruz9n
Z98xzJvXe5T5j7H+5g2U0XPNFWvldY3Q5jqj3Nqg43S3PgGMyNAbzD/x1ch+mNRRdSEQprvUNDZq
DClb0LHvzCrnvq1MOzEDX2BUq8WJt2v0/GMWP4pOrGv0SqIwycIgCFMCDxejy+pav8+BXdLHcC1k
hcGFL5WX34I7x64JIWeQMcnHexRfXGqAz6E6oA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
h1/KmDWmUuH0J4WzWPNy6MyUrJorCRh+4emESTIpt1Wa4mjPcR2Yfc1PJ35nnFGWVLbh/am0kWYG
uz2mLsI7uxQZzaVw2mALHl7xnuPZ5BBPldcGyuakH01uKIYENo1ajb72tHszh9zxNBBpVirEBG8F
Xe+SegjMKJotg0azRztfW/ahGAGSZu0xp5kCP8XOFVscw+36mCBmgXThaF0w9PDIr608p7M6Qnmu
Wcw0W6RD1t9YPJjQSNfme59oKluI6Cd+7dA2avwjzW7LIhCbq21x87CAx4iiyZp1Mf0bqBIOZD22
BPBYclWolWdc8ZLm7t5lakznVvMK6yD+bX9f9fjPXqbnRU3B1HllPX6Cw0hJHiRi/ZHccOwhxcGz
qwYooJAlXY0T0wuN5V2ZnSj+ApJvTSm0PV3sJqYA+xhb8tMDvgL/7ANwhqwCRPX2FV5TS238K7X1
wLhVwLWTxNzQz7fVzHwe0i1KB287efDf5dB/EAWaMMXFQfYue5Rd4FdOdB5hDVnRxO9tEg2oOTOt
JAVo62gTua9oPnFockrpBbQ9fqqkwh9nK4iMAzQMn64WCr0v7oxTZDv/+PMMdHUpGa9lDjR0Xvmo
QwXQvhJzUzJcSNTVi3A3SfLXcfFqepZPGZU0MAk7xn/7/W8OYpmawm3bPz40m5vDxhF1PQmyhOkb
xgq61yvvr1HguZDIzhGjdbk1AVPEy8lz6c9kfFacTWto5V285YBiOBtpW5nRNTuMR4JiDDp+UgNe
f828mkQSFVUdNuAuXfk9SPPFzTbuO95upphGNcQ8CMhkVBLwWKkfW0WzX+FjQ36okPrbf6ef5Yb1
HsCEm6af2lUaj8HSOWxXe2iu5/mk2JOveUZ9lN/rp3teyuntq9QRdfmgaabA4KKltHFG0Pqws11F
AI30MkV3nGsCrs1ubr2CZN7GsXtpHuaPdR6VDHKPU/PAAPA+6qCp7d7HKFgpZa0lLmoN9K9iIXtU
2ITrBGQzch0uLk2oUALC1xW3JwsOJc8hjikshRmbBFDGl5wrTYQmQMti0O/cegFiIMXSgBd5dvdI
0vMTGjeF27p8mTv49yEbE1DnfM+DCmZA0m2W+5rXd96F/r/tbgtZ8HxHEA6OHEnuEURllQbsV78G
RwjqVvKdrT3gQCobQV7wloe2QoD1aamEpoH62kJ9mMHEZjIgIx5oPBH1yVmjRgr69D3DScNBVHYD
zU83lko29uZe0n9RBCw31+aKq5iHdceTTl+uwsLzSadHcGbqUwwzWigU/MrjizgCrtZ3XqV4Hz0w
sf2ix8lT8g7vh9elZmpYCH766h5YruE19bxfTNdGC5eJiAJZljxgnnT5kSZpfAoE4F8Ic93tKUsX
4/wBBOtKv0R7ZuS6Glqbu/ETwH0SejKkexGPdDh/ifvQCVyOrU3TLT5DLVxvXKT4PjtUA7F5Bjfu
oORVhBPhrzKaWll26E1yXm24J3Wp6O/dUaIgd3zXIwVR1oMhgBOdi/xhkSqVI0LPAybZPQXfDGxs
obRlCNM78Jd8+HrDo5P+WhqD4xpKYOv7PflzDJoeOIxEdOh0DnxmshYvIb3gxytEAPOhLhh38A9p
KhCmtdvrtIulgUsx9j7RhtiUkVKHVyhi1RaJVWX7kPnIJpim3IDw/owrvdjhOBtZxeDmPLiXVdnT
WAjy7DNnTrWSxF9gqKNeKN/rfIc330WnX7KElX0h7YTn/GjoE971X1ESqaSU1UCAOMEnMjwV5F/6
hU9LS4MFUt3nIsMJ/Pi0Cg3d3bOJGMDNqCysw/KpnR/fehoOMGmJKPWwXzW4xX3edJl3wm9WHlUP
Adq9f71MWkqowXYt/b0l1XY6vGisD2lD2/hVDQ5z9UgbXkxELvZilSpUnMDyq/i9YmzNsvA5WtBT
IRmKHL0N5BTPE3nD1nx2XJVNgsP0j+LKf+zOr2+/slYqFYOihwt4jm3mJ+1Q0BePPpeHz6F6uyjQ
mqAAW1bXyi45IvoSFPOTdfNr19p6t+JThRjGyKzyZfoeHSbOaoaFnYd8kQJt6/jj7Md0gsDfZLWH
nRxGVscy6RttFquaLVvpAiTu545wCNLpBMoID3Z6nGIl0ob1fSfXMkONBuafNuzZ8ROgxQDwfxd/
r7SSxrUzyr+JjaZth7vcmpuAiwkq1T7lArXh/t9xtdq3oOLSl8ofst4CYBE1wCigKYoCyG1+avZn
pNiTod8JGu1IjT+WAV96IaYgrYTs82bVo9F+TZJ5kkgMMoZi6X+2ooOF9Z0GLiYnsUCpQ7NK3PeT
BCvkqlFprv98SoZXb7HNAGTWNe6wVZ6O3ycsDjCeWOHhcwgaQPnCfUrLQ7srcdipPIJIuh6C5EnK
WO8PdtveOCXqMARMtqj9RtVgIFa0sU/cWcc0BrJ57ZiuyYS8CnkB7OacMvfMSxsCGWOGtVnW2vd6
LPvMbIy8cQqyTQoM5hOTDX36X8RmNVyxH9fLmoml/YnxmmFpFJiGX0F2DjkC/7VwBOCxbgsx5KV4
v0uN/ARiA4j6/Yx92J9c7BUKouAqw3mgaHVLM4OupGye7EfDpQa3WhyBuD/p4MGpE6V0wHu7KnKi
MzdpYavu2nB3vULzqF1nFIipRQm3Rc+o7uTqCon0OcLaNYWB6tg28/Yyaifeugv1n+6HhO92pzek
dv0YthFaONKpjcee1O6NYKtwt221d5KhZCZSxIOWC8IogUulkFzXUtFrJgaB+J9yxRTXBZqT39ap
7kLY3SeZCzL6vUrKXe9MQuonLZXI5mpVEDeye1KIgCFWjyiCecujodGDqSEhMXkiArgKPobqtgYm
sCXeNjWXnYk6jMKVvjxLAi890x47tmzqF/fcv7YNwMPuq/yYmWihJdMHvHp6r334rcLJY6gY8aAu
pwwa94/hi9/clAuFIVnNC+dkFOINubA99huIowFEw9oO6A+U0C9TIeVxN3E9xf6IYCiZO0IKhGGy
CgREEtTwL2hH8JcaKgorWj88JRhCSvVYBWRsc78OTWp0vzDwTowswhaC9v60FLoVJX6Pc8lvYw1s
+9S+QcUY6JPJU0AomjPWF+0UPK5qDiaFn0ZQAb4Awusvnwg+jhdDIEISEbKizahaL4ktBL3VPlH/
JyYdukLWT6IExSASCqsgfiCqsidGQshDc8+Zg3EJZ7hvDRWYv/Trl3Rqrpf57EXYbL+v0B7sNRoM
Q1+F1jNKZhl6OHzbLK1ZS3p5m/TwyLM3ue4FyWVfrG0UaltwbtRkiamYUz7aEd58o+k5DS9NVeDt
RK6A2btp0xGYGjbA7jFkSh58GeaMq0JDQdNqa3AGgYFO+gzG4sKUKycQACKVxb3WWAbTO5BOWBOA
2/pvOu0bAb9DEOnuyYQXpnh10wmYL5ShWeTAjLr2nxrt4UDA6OVmHnl7Lr5wsl6FFb18mTX3nCn+
RbvGWlXxoCBurWXBcQycPPVaL8wXzKLy/eFdJnJCOBgzO5Tigfda3Ij4sQRVGWlhVE6gmBKr3Y7D
tk9YC4HO7shT/LV+GL821JfcGfGt++faNKrSlttbQJ3DD9OSmTsiDqnK42cyI8vMu8RzeObSN85E
2sZBmrRkT7Yw9gHbbqlOtgZmgM5qJxH+Y3buDo0GuCBsc9acvztVvi+yESogwJxzBw6R3VkABGN+
pGNB3Q7DMzLmjRxfgsXq38kv7ZxyTFRrfABmn94vjIp4//hQpdOCJe8uNPn1UjGMpDDMQhpHgMyi
Y6OPB/AtZZ4DdTpWJx2GNdiF8ftRGmu9EKfnHIxK/FLCZVHdJzgcyWuJHcitrprBCdzYczZzuY25
Da2rHtAh9xyj7Lm03VjfAPu+3V8N0PwqdzG9Z9ervPG1mRfZ2Bk59VTNC0l8eJpY563hTnOc4v9E
fXtYhrQdbADejKI/lBI3Fcvr/+PO3awrCSPWOH7iShwkKNsuTg0+r6C6LuXwjTYV4/v1CrY1lDdy
QDB+5NssxvPtTZAktXs1t5UkV1naDHTEgYJyVv0hO0h87tMIJSmE3waEhz9iG1f+AsucazfjPcgF
wub/sge8ObX48BO0+hc+vO5i6jnUfADqwinmyp/21kWUEr3B+4s5bxNGVvVnQw62G2TPTqrYwESZ
hNr7PgvLptqT8YrrBs/CPEv/ZGDq46iOOmW4+JKooIQGtsdycP5COHPN7WH2JzNOjHVTrnlwlk8s
qGzqmCivN525ZpBTz6pSf+PDE0hd3BZnWs7ttej30TvpkLM4tk2RsOCgVNn+9jZdi5HAxZbpq5qw
IsQTeJnjBZb4cFB/ZyYNVOb4/7b+eSfhZtZCzg3/F/xLxL5z7NLweYHYEhhsmdH6gxRXceHrWdKo
B0owGrk9FruiyWtvZnBLPEmTadQoM57/Kir1DLw3sRR0BpVl5iCuwIop1zzFvTKRAKyPcp6+mdsA
XjUUdhRPrb1PZmj1lEpOCMdejkrSpmzaGgqj0TO7UEv/Q54KhVWRy/1mh4+pAicDcudYNVFn4WLW
R6AuVkn3Hk+6N/SbbGvKdSByrCHNfQiINAa/N9s1H5Q76IGwd5ISr/6siJmilpgn7R/jyuwv2idf
8r//A8yIpz+3UCfJLYqi8Xuf2auMWxE/MqhwhasdQhduEoSSPf39buqLAkecjFM2IWrsg75OFrBk
2ZtZDS2wtJa2ykraSGZLDlP1U0yGiBUxBvzpl6N3W7IqsAzJ80skgjV1XbuVKUkNZ5LFESDIOo+q
mzfERpRGdqLqUwl5tvA3YvpOTujTh6it7qmaPHeUA79eAZ7h2Gj8Lvs11/2ncYgv+PlWt4OEbyF1
3NZAPb48EQ49TiREY7DQnQmzTWbuJx+AY1IIkwVlhNW0ysHS9PAQiOvWHOBOy5uwaaX4OVCV9mat
aPTpTgoWIxTimS+bMq75R+BcOJ0AQGVwN234cWbhcIreQeaP98fgzyARHVgQ1uiGRCwi+cG2mFlm
CdfOsDJUwjpi8BYMWsHji3sO/KmrGgEyJmejN9AlIc7ctdDvBJrm/t3BplixuXzdWkgxS0VtKHP9
dHeJW0Cqcg34s8f7Sxh5H8CMzsdtqj+n0xFEHoMJc1pi9bx6X3daHIwj+RuCBhU19vbGUMGrY76z
ppuESGfeymAJN+lhvaLRYJ1ThjbUE3N2bUzvtRO2wz/t+KyoKNChmHJHjKgd4s+LhuBkDBSOso/M
D0p0JlMDJempSRu1iMksQVtBsW4caGBLVcgiD74sc+0XUcsH2xDPEgPz5vVML358hgaXJ9HeEhrL
DCAZFbfxKerUsrZe5zM4yGMX3Dwmf548yZMgzOT0KQs/UngMLIN9nKwNM9wEKReavT75XUOMdil1
jiDVPgalZKA0BkHNi60RemZwW8y/4TgVp1xHqtSSSODxu87odaJUklATtURhu+42dUw5RhFgdhxa
7RpQ8yoyqjKw0olAFl1IFw9M12Jk99edxGjVFe9b55QxgPBF9OLQyQOjNHhRmLzDE5LAQPRJUa1q
1ujluwPa+87hhpF0A1EAwW+DQFXvjeHcKfZo9QSdFLTC4XdAPhUZTLdEBwO15Pzt81JM9Jbw3C3z
GAzaZHTAD1x5m7GT7kEqKnTFN6fYH6UnxZaU+LqY/VIxXkYjrzRrsg72PLVf/HoSqA0uSqDnaeCy
KVXK8ze8T8uQvq7WxYaIZd+LwjTIOc7C8v/VF2fPIMIP8luOxjLoi8mlbqWT3GO5ztf0yRyO+Rk9
4hbIv834IDLJCcYSYlmjBr1yVSU0aC6+xotZTY5WplscB9tKZmgh8sD24i9B3HIrVJi0S7W4W1LJ
2hNW3rWvAKFFHdswrL3E6Q8UsKmYT3KTjPc25TIItzhbu+XJGsVdggXhMYc/zvllAezoceUqS87p
Aak2ziLYpvvB9ezq5GQ+1l8S2jfannlj4mOYXXkLvmBSQV4BcqpLYInhZv4ABY9dEalqrd0hEArv
0abzTNkIwBgBdkub1nsl1j6HgSFtzaSIhGA+Fl+JTGxKOKiTGiHBkM1UOWG4X32Gbe61peG96Vp4
elSGyhI48Gu8BwEhzS59U2mQWj69vjtUghKRgdzNVbv9e8WpMpAvyAtGa+mitdsHlCfRi/89qk4d
W+CaQ1HWc9YXg3WODZjL2wNN7Ju435fZLTHanzHye1B8rO6VEMY8V0PkZAia3RhmKzyJmKlwKsdF
3NHvyep4Q6hoGepPgJycOrdkia7p6l7gwuHc3FSXMO9l1VoK4nVz+woY5yEbP7t5ga1R9ccJqdc0
ozurho8MeCy+k3J40+ylWF4Cl8P7EweUB3WDT0L1vGcx+m8xd6n1oN6C6IA7eMjny2nfLyR+Q/VQ
SxrNsraehmDe4HIB5pUbdORVcj5HwQha+L6F+hsXqslITf1+ZbThSPr1DLgILlWvluHPp/NLSFMQ
JLFuFvtcMmN0/tHLGQKkhAG0p4CpWjEeUBXHfKQThCl1VGX+Qq6jhpago+7oXRn608BDSH+jc2OJ
2f2EX9qBCTUbxHCEApfK3fpQgF+0Wjb2opKSfN0vVZihMGG3OM5HDGiBXirAF/Qgq5zupgb9eBjz
XPbHTffFefzArZ/6tEU2aZ/vbJHyYIYdtlWINFTE+oxvPosVOPU0TcgKGBP0En1G/rXSQqFRXjEB
T6IXkMN85afnWL9elLfhWDBQZGtdtWNDcP8+z/Nt4Vlu9SKCUjM7kUlxO/jRvgG5muoJ/o+fZHQb
xdlVPnsr4jklhJezILJGK78gXmUshPZNp1E71BnStkXCVIwZ31PvAv6afO05VYNs/0hwdWs6B0h4
UAqYns5XfZB5M+aeGCegCdpnlCHbMkq1Jchj18/fMLDGclTszJF5kkztkf6kvywm74oRCsdXxIYk
qcbtgf24++13NoM1Pe+zDSuXEQa3PUdtsvG9Rc5sL1ED4LUfz33EzaESlEKNVTkYzy9KLKWnWQTq
EwOBwxHxmki869oPZZAsh1hfHvJvV8hC5AjWlqEwA1m/T5VPoCLLppqKCSgJ80no31CaD+UJ8nGh
LxvJHbu35n2U1fbwEwOup7CDb3MFtb5pKi1QCjzdDSOvBI9Di2TFUT6BciCoWCJWwi6f6fp0WzAY
HgVQUPe2AUsVQqz2LtsFk6+oHV6+agJgOlmVJEc04X1jaKiRyAYluSQfW8mtRrQQV1JO7SDciL+s
cbccxnL6pDKPBAUAedQIXLf5FNDUXnFwEixa6pIkm1uuOhDmSfyGicx4us6whIoN0jmDl7ZTUb8U
o+yJdQdHMvw7NBLnNYyHL5RHLyN3tK3AkIQdVe4ntR3lizxIukkV403bxtlRkx+9rXZ3Kn9Qvgzu
LX2AZzeLYzE+rsHh6GjEgo/oDTvtynOVcKkGro2bhoBTV4MpWObPq8BC6wJBFPSR7FEDRRZAESaA
m/mKSqeCPxuT+qj6nnOdWgiWbduTFKkhHQ2IuBgDHn+b5L/ZUGp9gysKtzxPw0QYOzKCqGcjeo9G
5Yz8VP9dueOhK9M9OGCJw1sZvUIouHjJFBoR5Qvmcj6FozZYcb3HWJgf+S5wdyRm0lHGxoVtvaZN
UnrhnI7ME81bmwgKsTgdPwFEsTjxGHGljZkmJDjCfOXKLtcoc4N5upzeaFv0fu+z4pj0+volFvkU
v09/nx7u1+cE3nrin5VemfAl5OAS3q82K7dnO+CGIp9bBdNwLSorEts1fpEYjziJB/KGsgioVNhp
g2B1f+O7GF2uhjIKpiYgljTzboTI4hhME5wQV7Yaju79TefoBCaK5IDtPLBejRMrrVqiX8mRMyar
iU/LHat1TLGrR3wUvBq6i6HhCcnN2lHwwayNbk6qnM3mWdPbBe0LYu7l77F3sua2TVomfrqhl+rq
iSq38xrijwkEL3X3H1/wf/936lguCoRqtmJHxsUdkRUMkFyZ4KStKIEYVjoWLX6+no2hwVxsZ+gC
mgYku/W4BK1AIHKpqh/k+TdjDzA1V+cbZOSzDWzj24DjSVAntogRu0NLP5LlV9uAvpL/1Myjli9a
/CbBkvvFPtwdDlkqFA7aI+9BFzCd7oKfByy4uHQmc8EIOBRB0wxJd5P64pVDvUMYfHNszsLtW91b
6s3WwYBjdRe3XBUTRN6O6FYwydfcqmXtzU4Q4IWXfl2vkvRExJyp/T2trfFbp7xoUKErK8jo6OLd
Iu37QFORBx+9g5seqZNVQJSptyVFGt11owZmdIJLPvZ/qNBDRaFBllh97wfmxlgIpA094Ji26r2U
8V9fIJBhFFl0iomdyoljio23CCUV7E4PDOX0HIO/a0eaho3FvYZmn7zhRTjSRoBrbuYx6agnu3ZZ
Lhus6caCJezkCZKM0tqIN2Luz3kDeA7lWFq3/JhPAVy6OE0pUTvq3xF1efNjycThlunMvMGemoE1
Um8QcrSjMuz0yYvdQTyUpRLw1JhBhTwaEYCkQ9VA/E+OUY9iQpH84fTXrnyH5t1pTXoqxPa20u3n
Ag/e6D8vYoFknULbChN8vbISFiGYCx4aFGcQF95DuxanE8MQ7MuZyZpI2h9rTksj1uQ4IsVLQSyL
fjUkmfk5NbLN60DqOSCZZBu/xa28V66YXsK43nroTQAOxUYZE5ezuP6CKjAeigP41hz0/QfpMN7v
2k4a9k3RMSzUP9D7aAI/MbqrHeKIkDb0TGZ/Cd5wNGe5BRxJinBSJ6DF5N7IIo/ICMQd6FWoItfD
H985ir/YMqxFDl0/sAHu1G7uvXJRIy/UZ4m+5cbrO0i5Ka7c2JRMMOnU3q5POn/1vM0L90eXEbTU
SX+OV6ywpYKgdyFfSHfZdYH88OovYWtDXtClF8ui0TXmcv4jJy8s3SapAIXqmjUH2bVCrGf6PKO4
czYfl3qGsE6fM/Y8h3fPsxRbrWLLYGgO/UqAHKMphwMxnOx1vgrj9+oHuOT3NZeLYCRYds01Wu2c
2bYQ9MLMPxs0rOQmu1itByYT6SQhV+Dot8oeLI+UJS4tW5yVsv4Dzb3aWzk2fH7e9TglUX3GRxTs
FctIqeGG9KuYB/8Iun3ldRLgjJ4CY1U+76Ft/YUrTuLunJIzA9D2+Zv9qLpUYQm8qV6bQXATDrEf
RtnmohG9qgCeLSc/CGlrvTuKIAuxAHIeYuhi8gjwm+cuCewjfdv96zmWe5iDIzoxlHBMhDvPgs7/
T+FeIZ/qMgs8tT93XRYaTanL5rINzfnlKPQikdHWU/3U+j+cfh3u6USQwggdosyS3w5zUzVChv+Q
ufb6prvRArDAspi6dlNjQtbfQ/Q9EfJxZ9ygNS9ie2SiScE9JzLSqxXo/P3X+XSZ/jOMjRsD5k9V
pnJvMVBMdjEaDT89bp0YppvKT2kofTWTQzQ0dFTtHotyRJdT5hO4Vmt0qM6zf9mzqa3ofv0jNy/v
9tfJ56JcDycTWhhjYArLtKan19mnrd+8CBB7xkhNSTJkyfF05WzDzyN3w8kjKxziHsCNa4NACd7y
ZR/Ohw6PwxNzkyc5n54lghmffTu3n8QfjxQTRh4vJb7okiaVv33dOru2TcLI1Hg8yvpxtdjKETeb
hqClea5YOLWWfE94/fRnjYvkeubLpPVSqyKYKeCAv4lPADzv/XxUVSEBAPQVo/kvlojt3A21zfPR
ss6hTmT/EPyN/pEiHHUdj065UcNNUELQf6dwviDwSokCPYNhB30NZaRoDaiSTRYIamG2rhdawNud
2wAmy8hx4JXiaMAvwttRPE68/CMcjGyGP6FVyaYQeqgSJe2L/GG5LG6a0UhifQIZVanOFQviJx/e
osYJFVTMYWL45TqPRNJRiRZx9OzW3wUsN4Ptxvhe5ZHdgg7kiDWbUf93DEg1hZH8NaBIJNnsmgho
nzpM6S+JyVcazyKL0RfFBMa074ZnCMRNFjQjfI7T8lf+flXWFtCYv+NH5tDA2CAdJaFePwn//iAQ
5jkzTW2VNNFgOiKBhY9vJeuXw5rtFwpWOfUcGa69aefaWULCyohBNxb64U8Uw3WGsJW6AikrFPpg
iyUtlTy/ehgw1af4RpWGboLhVbWMjCHfinMTJfakt0++lxuCn5stupvIb3WqLvTLiN5Xr/oYVVS6
hw2wc59pumww+tKsiemabRTd5PAyavpjRnEGh8XWOM9kwHTBeYYwwZvhcqBeVaQqF0Zh7SHewddI
u+TejGAW0shHCXsk3YlTT7Y71F3G8snSsI/KOCZUebTnDtLlRsSNfr3RPYYQ6VNr75Utw10gbrZa
fHAdGitdCDq+6G7rrRGOyOaeFLhXstqCZ0r4UWMlOPrwK7Tmyre0gmh2FPL4RrFddB6XRcnd32t/
O1OCsphiqxW15KoJv9KwcS6Fj3VNSC8vjuspTvA+6cizwyqQGQJP9Sd3XAtQwJLfru0Vz1zoisoB
/mJYiPDU6xpVHMxqT+EmCpGsH2f9vZdrKPmxPZOY8s9jiNUdI2RHgs8hY39cFZcwCsaP4f6j3OBB
wTIav5hhmhXLFNF/l4vCDJWTnx1MYDKCN3o8VZCkbco8krYRGIpE/RbNx6tp0YYyvam4pR9gHU8B
ZnTUeP3KGrupRLK/0A1MagbWKVXq+gkJAeVmrmmOPR4XDYSufDNDqLpy5HXQumVdGbC2L0AhTg6O
6V2dCuVqdyh+sDQ2hrY4kdxg2jgKlh/fJ7XyNb15cA9eNqyMvmL+Nr3tHYWVTMHJyHfhg6FJ4t+u
J4OaxiUulkK7MrBhI9CBvIOgJQ/2q5FT63y0fbvb3mpOGz6orjDHiyf2CvfGrH2fynkH/VkHaa5g
yZvmA6Bj4XFuQTHvh9wYXv3+k3u3a/yj/7JimyU+hwotEuBgSlVTyFfQ0n0Ug/WHpF/lVFdGAAvu
ML6jPGlRIdWWI3CUIvAs0pMUVjtcsorh2kYxrA31JNP6i6R1gezj8MG0hgrv6A+TYvPNFvyIvA8A
G4j40yM9Eq4jOIkUMkJu0q30oesU6ORuKQsf445oX9TnTOYTcJ0IgHVGFsmhXvVFim/mWef2Ad4H
Oo2/Y6Elcszh+OZhYlu1lYks+E9V0qD3x1Zfo0IcXhnShHyf3rSCoQVUIlDjVHlUdtCZVE6Fj61I
rNoVT/fanFBVLiMUZcdfFbV0L7RdO3zb6CdXPtFIyw07IKZXRfFD1OvUyzoDRbwzvoh2i56Yi1Oh
n2t+VdGnsxRpU8yLnxg+acdko4UVPrwoXmQMmAeWowPjRRfJHsSjWQeOZCMW8tCf7FCxocZfZrEd
M7wG3C+lgiQMr0M7SNPktkY/A+m1Nspt/+5/wIb2nQuc+EP6hYxQ0JEsGgj+dR9qTrYFJ8WNLI7M
8B/pu7hqpllEITh45reh2L4iHkCaHVFJmiJ8x2OY9JvPV8LlQzNB6FsDITYejAJk4p2s3e2o4/Xn
jI8l4bu8OmrYrYaiVsDtfwpx1YSpKW4rwr7X15TkNWmuiLNThDz07dampDyTgFtWpTYODAaxjtaZ
K+VrhEW1v+AAyldGWZlYYZ8NsRNU0adKs2AnLaa/Id5N3SzNcOagHli0JTJfNU1f7zFzjqn/FcAd
UJO3pl87JCkP2o6VFOUUb5vhsZdF9aW4VqSPSonDYx2fLLOlKmjLgmJB+F4uaUxza8ICelpSkNiq
vpTi5snvU38v2Y+ejo3XTiJvu9uEL33T3I7VzFtD47kThwVLAPzPFiXn/CI3c7lfasC8PAbwPQhE
0xkNo+OeDWHx94SE+DXBM4UlYsDbAuRrT73i0S/TkKsAYbb7KMHZ8uUNJFXBHHMjkBd9YS6dGlHb
A+J+jcaF8mqKTHM59B+bep819IzQNS8okP3gsHkjfJfhtDNWOqMny+YUO2XJf/5SAc/VI+ROiKG3
F5srapIbVAXOYd2sEdpNKeZn5hW4NGuHrsQrXUS32zTmQpyJT1kcHcBgdNZOWhhPYjsPLW2oLOgi
9hhwO4uRORg+q223kPKeac+HuJ4FcuCrG5IOmqi64dItb1nrudTZ42zc7OnxoCuPFuYt1UvFPTVv
SD/TR6wu7fAzmZwSrj/G3vxY+86ljrKODnRuAWxxiTcRF08DYHm/JEN4kqVkisrEsZI2X+4jYCXG
qpZZVVQqgHRsErz/5yJLnFHJpR4jCaUUgAiKvwTGNMwjvm81CyS/XMf7DP14F4vKnJpzFpp2ZiLu
loF/ABkLiNIjuxxjXdbda0putmcRpM0/7WQwbsls3oO92nuqanmNS3eiyJ19+vCEch95YxTaL5Q/
6eBRyM50R/EQuiZQDA0mmbLjit47T6irmpbjQU4c9sTd/+2DCneZw58XCovmqYadfHlEEEqp/iZQ
Xj9xhTHii7r0sXrWFoq+G7QDL0iMnSEQcNGfcJcxNqFC0vfMCuoj2fO9f78itWyXXjVg/oSnwtiw
GhBK//X/XRK9ZHXALtCqSZxRiIG/BLJpAmca1Wzhlu78Kk0HmeSNgwmdZjORcVK73SBF3SWtVeVo
Q/XBkB7tePxw1pT0BZN7UFzODesvk5Jz92blpkBBTs6xk4Y7D8kaWndSWgMEbJ2EMkt6Nu4kTjYf
S0KirzqNt4kdCZLFyf28MxHDRyIf7qELsToZ7+AJb5KfRRoZNZNXfwbXK9JsJE0tBSLs2E04mEJD
DzZ8BonYyJL7RrWfvK11baxSLqj3Lnc1oTJj76bSdnKEnFzaJiX93lzrW+OR9v2Sb1NQmTNG44zr
w8cH+B9tqndJWf1jcIV6O6wyOLz2+GPCJ3I86XOFVkY8vL6aGhU7BhSldzA50wg8+cP5WoifORFl
lYhDhbvTIWH1OVnbs98bOej1AMnBX0dofrHf777xx1kWu5zfhE4VlI1HdEu/g6ASQAEEGnxL3bGo
QP/8XTEvrPjyozsD8Q+/iSc/tzzOQ/zWz+Yq+8tYJnbppfM+Ypf3yAJwfn2rsMjOXg/sS8YKIHD1
0mz4hRLEr7Kt+1AfGfcAq0QjhRxK27WxeroQI/YLTSeukNy3fwYe4TE5ovQ3l5GXEW92G2HhuZs8
D8ihAuFHksaYaZ7w53LiPJnMEXx8mIbue2FkjJgTRdFkZzvFPadvRZ1qkDnuIyq0DuBszPqpFsWj
wlsl7wVRNC96VSNVN4SdQQefrVsUz9Hy+xiDb7ksKtlLDAZDwgV0e0Uy5YdgizZ5qCWKxGQB3U3m
5ljnz7DBCtrXREB8WLdizZ38K6gqSLXOJUf9gnDdxu+TvSbIFezk71eZLsaUPHzTEDxqdrVZ594E
+iM5u2SG60rM909CVD7d9qfHlB5tESbJqE6uIGz6estbyrlVO7vbDBILWihERDRErI81k4O1ORJc
w871mORsOLcX4TykxzTKG9/yTPM0FJDMITbxIIC/Vl5bGaKXHNgoj5zValc8UZeff+sVSPHWJd7y
K8k3gPl+dKqDzSkUMqx6KPzeIuwqJnNBHxLbo9NjLyVflPlnReD2pRQT0HWjSDjnyh+YwvUYTjc4
5MvWLzGAKrO3H5uUYN8AAg+x81qk6io3XeCsZw9e/edmb08ec3KthAKBTa5nhThso/e97cupEggw
7s4WUzaVcBS0q5LN4IokuTHf4oenK3xYXBL64kK3XU/LM+VHCs80rp1tX3f5O3Ud2lMxReZ2vP0v
pirW64rEMp8lsZWy2EPzD2A3O6/lPXKsGUFoum9MKkwxY6BxwfRcmKSB4qLjocqunwRN/T5AZkT3
wFqHM7XIT16kcE+PzCyp4dUu7/e/Cl65Nz9eoH6hggvt3arRJbnPMUEoj2owBOOlrixhylRKdUTz
gr1beM1DdBNdN8g91iFjh01UsxdHHyAYVqaxRvckfPiesUUyW+QojWXYIi8SD3nVgx4eaJI28vKE
0MWJGz4PGMzryXrHRdOM5L2mT6W1prNXDxq1uw43e0HHv1drYwgh3sQ71zaZn6+NZvyyjbvBqr8h
+tdaLwFJWuh7FN80blcnmuvYvRmUhJ6tn0U1s7Ae30YBUwbJL/vyUCFA3pM7g2WwX87EMBE4GmG0
nDgCYc5Ec0P72TyalXrjakCJr5bHsSh27CHfGMAoEerlGPDM1HuDFaZ3Vo0yG9Z5jBSJMFGpgRix
BeWzscpQMtT7E66PEHmZkY/cW7Y/QQ+73YnnXJLDmHyMLVuaU7CHbX3aQbyW+efhUoh6D8mJwBSU
jhy9KO3s3k/V/jXti5TPZw6Yj4S2qAK7f1bYZVI7uCdLmWSXYnRswvSy0cC8ylxQtEnBjircM0R+
11q/XG9lR47QaDX+1IKHW5e+8boB4A7sfwyfIYWpp6X4BXgapsm5mKeUmhc9wEVh1jQcrATtYgH8
/ZmcIW0cTNIX1JmHSw2o8NwFWMJ9WytmfAYfbg+VOwQs0kQapQqNXSi/tT624lvIns3ryDarhZx9
no6a3ogRh40r4rLfCEdWEZdBzLQJ0xptz/t99MfobUdoqBxGoz7G84D+a6KqEeXpDMQKoezWjKxx
q9Tt+xQeZIf+xvjn5bS7sBPvK13M/psadC4dwyzKUn0EsLwTkEho1shBQEfPtYhqemrAqaZBJ6Yt
wT7XI9K+cbvfMw5DNbGgj2La6W2HmaEJr4XjEi5Z1BgOu+qenjJ19DVwBKcjP0cjcJJy7zkBl2xK
bPAcB+gjDILePvG2S2quQ0gAwA2fao5C8OyorJP9FFDbV6qlZ+LGggJR/DF2kau+LLq3WhRCwGGc
CoVLSebL5OR4cLPi/A0WxM7zmMRKVcGQ9tyGflyCP8q9CazBaQPs5aZOFOGQnqjgpuFeu5wqK8HI
N0QT1qm/4G6YrdhSQi1q7LBcTaHw/mgV9n6jckdJTHDudq0bke8xMXn882l0tlhUGTD9Kv7p9Tk9
COvVEtBGdfAzcNIy/RTBmfXgVTH7+1DbuIua3QP1XQ6Lc4H4Wr5rEtCQXJDipGEXnQETc4VJc7XM
mWpv5w8YCpMuJ/tpt9/xIeEfZU7wAYTn9aZCrgttk6zm7szc0OPIM9XM5uzT0LqY5xmm4LGlSc78
z18JC64KBpSL1KjazCwVudLVqRvVA5/4N0iexb938OQvOGUrQNVooaUpr1cTbNEW/ayXzccnB6PX
FMLMahik0ScpMGZlX3/OVIIn02GBJLzK/grDB2+9LbtEdvADdWnV+kGk/mRI1jM1mEEp7Zf+fXJH
6dGCevCstiF1y72Vxb/7OQHoetyt9Bk8fD2j/APfzoICV4SPzdouurEdbeN6QtmCilz6nTiW5Wy+
Ttlpqxc2QNDrgJT4zhS0THtizu7epZFUzFLvk7KGN9QuKJ8I0bdt8ovcU7uJU0DTHMgS1bVTdzjn
xqhj7Rs8Sd5AoLbKrctmiVrAMj5DSyJO1RBp+Cj0FCWlGDiZJqh/hE3F+Qjn5KswluIA4lxkLwZQ
Ur50rx+1J/7HLBpljjCELknc7bzAjhrOW37zTvaSyNBPBOigi11X1QfcMxzkGn8692ID5viRoNB6
0+V7ZhTMQR8DQmyXA5q8EWCAAweckk1/0cVcJ1ChwfdGMbNNG/ECIFyCY0HYy3/3tNg8qBBPgLCO
qjBR4BEEpbmNvjCfZK43XEimjgDFhexz8aUoP2/LZFJO67mMBxpsmuBtpsmuN5K2bVVoKRrqGvuu
Cbb9laMK07fAQQsLSFi75NoUgoZFsLwUkPoa4de2ghviaa5Y/cRyYQYIndZ+sVvrom0qeWLePFUR
F81TjimyPDaF2xfmtAtri1aInDExx0XLljAIMm8s8npRhLvew80YL9kt5Er5T5x6KTJkCV1sQy4s
8i8xlECMoyLUJs4uRYwDtAzyOhm8ccaZTyT0N717qa3i2iXkTbaQEuZBXsyZxpsg2pEWqTKRt3xA
VXsx0g3SY/actqhxgySSDKDUYVGGyvd+QUM/C1/iYAX0cTQnPDtjiL+MMXg8xUxdDg0XdEHlZlWt
V6+mMzwikW+1sSBoyvxwZR/RcTZf3BSdRrmbf59M7+dIms5mEjjZsKpkom46gEx54pfRGxICBYuh
Gw6sXJiOjVkKAu0AuuO+rQDu4MCm/9qDa3Fya7MxCmgvuWCHTerucxQkbJN+8bdaVmoJ2HqIDiRr
o780OiW02hZhgNvZ8kLNa3at5UMhTKLmB7Kf/hHLcHKRXL6JGnmM/U6PGkk6rzXYzHW3OMWn0QgE
+VR/g3BCLRYYSg5037ME9zWtTOaGfTouuP63vyTs9u0ZkmFDSvXNOXe5J5/I5YnFE8b8D/5pTNGR
5gBxRP4MYwDFEwuzbRGBxgGv4yt6YCwZQf7fPNKCPa+ajkjiSr4RZDUuKFMZOpLScoWA0pkXn9zq
rpSAd2WT/yCLshn66N/PcOPC2y43djVkx3JmD8MGVRyiOy7+cNrViZphh/+fIFq6lSPjvzSP1OXV
Ozhaid2yRUOKocw6SzpuRaGv3V4ceoy2I9IxwGDby9FhKKEVzdq5S6cN9U8rtSDh09TaxZMnSNd/
8268yLVkzLFBUhYhwVnFSZdlrsnBw475koA0W66+OxfCZ/x9osMqF3Tz4ZCHPRHEa/5ylx6tuWch
/0u+jFcb6pfG7S6lXXe8Nayb3RYDk3ngzKD4hNiFR4TdEOGQ9ps0QwW9+m3wEE39V3ca+W1cmAHj
FCJDt7gZ65CDaDQTvzQe
`protect end_protected
