��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�Ts���d*!�_�2L\����X���G���{���2��� �buw�2NfS���D|��݌��(�)s;���A{�Lݣ6��n���M�L�S�@���'w�a=�!�g�L-��\/�K�c�3_�hh��@���R`R�����f�̘e|���k�a;,�N#M%*���6�@�C��H��-�Q̲ĿE6fX�?,��tN֑C��$	[�c�Hza�,��Ծl��a.+}Jz7�53����m�Ii��3Y6e*�5�y,���ym%I��X��[�xH� ×��E��5��r����Y1�>+G�k�ߠ����P�Q�/�uʍ�����AxR zRŪZ��o6�U��Mw�����[ ����8���y߽>e0
PϜ;���h��8�pn����"��+ݪJ�������Z[!<�f׀o/��&��n:��-?XadHL��g���}�`�7꛵�֛bw#$���i����(�lY�Jr.���o*�Ǜ�h&���j3��V���e�\��ѫ�W��=�"�ʏlا����[�j�Ŀ��o�h������t����uj�Ł��!��uoI[N����I�k[;P:9j]w�
���a!Z�ȗ+��w 9�J\� Mj6��un�1P>���$� T=�8�M5���,P13e��5��a�v[g��$]��ca�TCr
�z=ܷ���R�\��_��~�8K��Z̜C�����0̡��Q3�e!�è�5:�-����� ���.oq��P{���]�;�B�Iz�g�@��� ��@�[|���{�k�L�D��߱�x<���>t��QaY�#k�@r�SQ�+��H¦���
>=�b�@��:�p��@N�+�~����(�g^�Hߧ�]��9�r������LK�� �ʳ���1S���jO^)�2Z� ��H"p3�U�Bk-w��=�hP�F��_#x��А�!�j���:;]�dwV�Kp��V�&�W�i��3����o����m���μҮ�_��|�"�ܓ��k���
N|J���lg/(�2%�F�F�g.�U
�W6骄�G \��}�>@��an��	OV��]�!���1��9��[��4��,����"�V�nb���AZ����'Sŧ�B��,���5;�'���?皟P_X��h�����j��)ѩE��VAY����*�.!��T���$_�����,�s7WD����ƶ��4C���=	�!i���c��F*��J��#T4'�w�+��t¬1��g�������u� }BĊQ���Y�Np���%�\��7>��)<T�]k9��q_�;���$�0$y�(��!����j�]ץD+�W�Y�s�Ԁ��K�<,�����Wc��_�\��}Q`E�����%#<x9cS��h'��x�`l���М�z`�G�!�n�|�*ܠ�k@��Җ�T��@�>�f+w/��SYlt?yI�s-/�B�'�"��A��m[���`��h�W�B1xA������-�F�T8��vL|I$�	 �h��\�X�Z6��p��KsG�St�3g�R�����']�EKɔ$�C����⸽�9~�Xכ��GŴ�0=��m��/ټ��PZ��h��M^�?E>�<��R��4w�}���d�i�h������237��O��g��~=��
e6�ôN�ZZѩ�-��Ap������ ��ظ�A�M��!I����7?�2����q���L%9x�0�E)�	̃���@�z�5H�z����~��VF�˿�BR�/DC�`�~~��pHb�dqR N��L��H��|��X=)�
����2�J�v�J�h/o��!�\掃E>��PD� ��}d�c���]�[���wSK5�ho��|�Ϫ�������N��������LH
���m�*�,	�{+K]s�]�k��}fF���qF���ךJa{`�������oZ����-���[3�`ק�^�M� E51�/m�����HR���2�G�B����)~|(A?�r,�����Rb�x�֪��%rA?o���o0�\1O7%�T���k� -�9��h���-�S�Nl.?�,�1߾Ĕ�4�Z͌��5OL�~��du�*�!�Tj��Dw۱i��4�D���s��k@g�z����L�?ќ9��~��S�W�C�[d@c>z�i�o�H�}�'y�,��n�Jh/A�C����ķ�������j-�Nc����f�M�m�Ϲ`ʔF��d���rG��Է��WA�t��sI���n�$�*���wwݞ�4Z\�ҏ�H�T:�[ �6�ܻ�ʵ�5|~np$ �K�Co�b�:����*Z�>��
Vt7t"����z~��1������a\��:
#�n��e0�Ne��U�g�3�9�'%6m�	��Xϡe��N�C��ك����\\`�|rR�
�z$�i�5TŐ� ��A1B���_����4-_�d:����~{�j�3�?�3�*�}�z5nf�K�x�:Y:���[��Fi�-�s���s�Ǌ'$=_�:G[h!7�q��L��"|}��1�v��S�����fq�\�BG,�!w>�¬��$�����t�f"�����M�1y�6v����g��ھ��>�ޕ�z�mCU4���G��U��9��H�sj�8�Sz���Մ�p�� [�ц� ���VZR�b@0!���"�,��Z��-z��������;=����]#�3�q�s��n]��^Xݙt%��z�{��14Dv�v�r����^���m�ޔ2�/ߙ���\We����0iE58�.���e����W��|��ђ�3!�t+oq�8x�2��{�D.!�1TLIt�҂d�q�x����0��[#�yҍX�d`��N�`���Y:��	����%V���1�CZ�x�+�~��b<IY�ʋ���Hs� n�<8�hk����(�r$�gUW� A�z8�Ola(���+|����>E����1+���w���č���tcA��g8$wT-s6:!���_Xǰ!5r��� �:�Yᣐ�<�;�OԶP2�b����#K�jjiz�=�lT:�.J+��I}Z����x;~)���["�E��?��$S�I������[
�������@��6�Ѿ��G�9���ß�JFYTuz����*ܙC@��56hO�k`�Mě�UG�J��[A�>��:����2�	8��"O�����t�7�8���������~�IIS�l2���y��rg
%�Z���V>:�D����I �VRn���0�~qy; &&~�,�܂��x&�2(�������4O�k��cx=l'���d��oR G&����%dEb��r3/�	��Po��+�3"J����M���?��}��C�ж�p����>"z�t0��\�\(���I� �0�O6�޳2�iKjQE�$�R�{H��Z�$�#@�뜖��ֽ���8�v�>�FTU�A& �F싚-|�w�ͮ3�L$6�p�V�#�;.�D}���i�l�X�>����n9�1�' ��h��FZ�(�mKM�,�a���\����i\�ЧX�$�'�Mg|��]5QcE���_�Jѹl���,6 )t�����ag��e�3h�8c�:����C$�r+l��i���㿟l�U��+#e�
�G���c���f�P*t��Տ��l� �@�i}#+� 1����6�ֲ��,r#�����E�
�b�(�(�B��V��+��
i}L�G������Jc��$�$�������!�DXד~ٍ�NۙҚ���S[[Gp0��nM���Z�%�*���]�T[��ю*j�u�G�Z�sb�7��p��m�8m��W�O�Cѩw��r���� ����2WB
l�zwMQ:[�ʍ� ��T�l�����Pu|f�������B�����\z���$2!��(H����d�p�Ɍ�IIJ`S�
�I�[	u�Ppdɉ�΄�q��5��?� v]�;9�h"�5]�M�FO%�Jm��Ջ������2J������y�d&wq�@�x,ԺQ�_%��O���w��sF����4�n �.����v�_��!\i����]��N���Z���3'�������b��^y�_b��߆f�Z����h����YY�2Q��=,�l�|���_�Q�V]C�?
�-�U���efU��.��c�fV���5���h�kh��JO�d��&{=u�o��S��ܚ�Z��>[ �\ȡ,����P?c(��Z���E��|�^}ʃL*�;H��	\��������C�~��Jog�_�G���dZ_z�I�P̄����	9/Q�� UV���l��k�Lw����NgV��t����[�}bKT~���No��x׌,SJ�����)E�������n�i2�d�KE�J)U?��JG���H)E�rk��z��Q;lڟ�No�pw�����]����X*��_?V:AW��Wѯ��g�b�΢i�	�;�KƧ��������w�pޙgƦ������Q�`
f�ͻ�Y��Eا�=n5EH~*�ql�۾�\e���|$�N�s���_:t�52���-M���OS	!bb�'��D�ݠCvn���!�;�a�Fu�����9Z��ׄ�56�N���^# �<0��T鑆?Jm(E"^�Q�����^���Ź*�S�L��.#W�d]�>@|��9�3�M����p=$���F������ՓL��a�9�F*)�ڬ��1�6@��E�?�w��C_G�n����|�vG���?��6�ml G+�4U�,�1�a���Z��d��Z��S�գ;ڵ���h�We��!�4�����6�R�Q�..SAh��q١y5}�����N�z�=�����<�ٟ�8�C��Y��!+h�3�o��
�+@�Gv����'�ߐ�v�K�w^q��~��{x9�Y�S�q������d.'�EB���m��q���f�d
t�����>�Xy6�)�	f�D!�$��FR�	gH�+���߀��uC��H����Gp�4�'m�,����ݐ/E�Lr�{S��~Ķ��?qtd��,�ƃ7Kw�4&e�;^Q�DޑU�	�ob�R:P�9�rǵO��f��]�ݿ�����D�.�u��MY~��i�����(��'��NI�J����Ի\�".����t,@t��;a�1R���������?Q����}���֥�	�"AnH	���Ҫ�S����%f]�q�6��~��9X�{;V6�x��L�kd`�����<j�����Rf�����奔7��fC�n�5uŚ��}}8-^9t�>$��#�\�4��� ��DM�:;�m`DJK,�Moɒ0���Љ �A�z����&���CR%��d�d:H �4��<z>��Y���r�n��J�4׼Hz�6��49L�L�Xy��%�����1�,A�\��X�e`ԫ�F���dum̍e�(����+�]Z�H~"�T����p)~҇�}��mg�cM7���?XU�N1��'�W� �${�`B���D����@�WjR7n��Z^�{-�w��!$��2��Ӆ�R��@c�*����0�p��>�����_�ѳ�@�5���c�\1�<��~Q�
�R[��P��G-����ܯi������ ��X`�cs�����<8�^BZe�5��,�N��g�4r�X�n�����(��=o:�^�X���a�f������+��-%�R;O��w�Ѥ�^W�1��]���߳�ȏ6E��M�vw��1~�����a"�%����D�O�
:ɬ2GJ6���C�͛�$��.��o��C��3p��I������7k��f<�ſ�zb"��6fRɐ�Wi�Ad��j���ť��qOf�N�����n�v"8���w��>�̘4�wmr ,��|c_E:�?�궆�c�I��Y�zF�����1��<�ֱu�c�#Y��������O���@>D��+����
)���|���`wE(�N[���.�����G.B^	53ك�8�̙X���gogB�m����/F���.�u@�!�Iii�"��n��#�:��Եv��y�+7�ڔ�3L�	/�V$&�Cv�Z�J-�v������*V:5@�<�k�`*�,�i��ķ�e�9�v��ۋ˥��?v��!����O=�+��Ӻ�`�'Z�n)u���o(����8&[[�
�$_�X�r��@[P%�{�F��$_Э�㍆ܴo�g^(��͍�s1���?��M�(z[��QR
�2�;�X���ER FM @�d�l���q��၊gq#�ڍR!&��o��4�k���{:�*��4Y�}<�GO	X�����i���̝?蓝���,����W���+�����q��7n4��}���+p���~���~ڪ�Zz�b%����v�Y�N뱃X)*�`������=R��(�y_QA�\��9s2.4�R�#��Խ�vdN��8�V`?��%��������zl�и���'��u�ԑ�0���:���/���CvI�����~luz�������B�X���6ϔ�-4�"��=ݷܒ�ͺk%���+u7 ���ݯ���o��U���w��3O�v�_�j��A1,�u �Y0t����J'�AA�8>\w��J/#W`��b�a;82FM�O�	:W��*G�6�=NA�z�xiɉ�C�l�y%��c�裨C��ޛ�}�E�L��r4�U� 8k�R��  �V�����>�1.b+��r�P��bݪ�߃�A�İ�.��;�����j�t���s�S��L�h��[���
��;X ��$�wF�ZFB{��Gۖ��pw�؃���_9�Yժ
qﮩ�]%��3��P�������2��!��~�/	��XFa)��O�x��G<3���3�D����@����Z-�sb���R����ͩ"dT3l�m�5�}���A��I����VP�+Q+R%����yr� l;� oՌ���9Eɢ���)�Sf�;�h/�N�ɹ�����~4�1P���Ɯ�A�jl��{����@+�k�F����~Ǫ
x���� ѣL��a�t.�HX>�4˥�$����דj�޽�!�Q)�f`A�mj�t�6�X�p���Z�5&��S��K� �j���>�- ��w��
~VB�����,rZOJ�I��r�o۰t���4Q:�^1���<w}���p�G,ՙ5ҥ��޵�!�d?9��2;ׇ���Q�#��C�w<�Z�뎮�}��Q,'�;y���W���n|Ȁ�R0�3
� s���	*TQ�����]o��/��\IĐW�P��N �~g��0]9#��y�jr��Y����(�u`SD�yd��A���D�]�/�rQJ�D�nyh)Ӏ���bgZ��R��`�����@bm���u�s��U�&��5)	i�2�0��L�k.�xS������nF����=�^��>S�m�I1��Nw"��<�ģo���L+�����V�U��*�W���떤��f��{I�ْ����V�#�����Z6$R�2^��ֿ�8WZ�[�H�.�
��{��ؙ%]�7��G�0�'�{����|��*�R��3�f����J���ry��
jC��ԛ�!筄0���Ma�\I�2��c~�_��9���kQ��WK{�H:����>Z�^U�1�~a9��x��s�S�[wAv����{ VDݾ�q��Y-��t������)�<\�_���Z�a�d���PN�VSc�`C�4$�%�g�5 �������OkԲ��fi�_֏?�[�fs#���h��`�_B��� ��P��Wz)������+qG`������E͋��z4�t��<���_��	�@
 K�LsM������?���@�����S�9O]�=k�aˍ�1���+���i��͞9�ap��=���C\6�[㑹v���R
�"-N�����ݏW$�~KE�Ҙr䢽\~�7
`4�yJ 3�F&-R�hUu�Ң��=d9�T�jpՇĭ������3�轘l҄pW#��.V##Y�t��U�}Q�lj���I>�� ��@|��j�B>�㠚��J��iZ҃�����A��ʋ����{#vs�2s������'����p!ֶk�G�9��O��>�\~�S��Y�5�D�-�#���=���`����%�Kk(G�� ����)$��p�1�OǷ�S�i3���y��|W>���s��r��i����d�BRs��Q1L���w�d#��1�������bb��n��1➊�Vʉ;�~�چ",�[A��+���O[�.�^e�����o�)M�K6���g�4�-Hc�&+������ *i���h����l,���~H��V���{�M�,�@R��P��QESQ�KM�ıU���l9�tIi�-A�JWp�	��}��X�2*�ə�(�g2�Yi��v�F��v%�̊ڙC`����cb3[گ��I��Tƞ|�\.�e,)_�nm���!�%6���C@�܉ئt�ؙ����x2�b�v�گo�Gesb��2��=&"n��bE_5Q��Ԋ�"ȳOz��&��� P«�}0�D�Q|V��J%ka(��P�tB`���]��@1x�R��7�3I��NÜ2��u�aS=	"�Ǉ�����.��u�d�ۄ��������K1?����c���,5�<���G��/���\_�)wi�v$w6d�,�r���z�6鈗�q��F�ף+3CX[^u��hmݫ�Qg �u��3N�:�ěx"�S̝�`$�r(ć��f�S' Eں%n��6]�]M�)�d�:b<�Ը�Ǒ-J�^A���G��*~y�܌�b̔aY@�N!�B2Y�[�Z���N�7�}��8���N�c��x$`t��D�C.�\50Fb���bT�6�C՚�%(�R.�C`RJ�����*��D��t�g�z4vAI��5�������w�e���W������&4���y�u�u�Gٍ�H4b�	�����G�?h�pq-����6c�l��y�=��%e�&�ܔ��N/`��*���1_zƤf^��4,�Ɏ� �^��Tҳ�_o�7���KR��(��K��|ӰR�(���pZ�i�1C�Dl�\��gT�r\��xzc�������^~�[đ����[��Xf�Ł�a����Y���6����&o(c�_��鐜X�a&�OQuO�ϸ��>��y��<�+��ʝ�.GI�x�x���3PCub���()]\�<�(ϊ�)��s/�%�*����Gz�������J���4�� ��B�	]��eR������"��ΰ��%!�D��Ʃ�(�>�4:,j��h�FOt�&�o��U"3Lh�3:h��ӆ�=�+�(��e��2n\�[]"9d�Mc%��,j�]�|v�!�G�>����w�2&�~>��O����QP�s}����`tx�6��X�7R��]�a��ć�3����{K�i�������\�3�e6B�L�6�µ@^�I|C�Ϳi^���w��d��0QI�}"��<T��R��T��(4z�D8��Sk9ݾqf��U��@�*Q�l?|��~�������!%$��J���P��Ϭ��;lZAH-|����y��%���#Yꓠ0N�NVE�EE�-��m�����w�������ͧ�-RFq��aH�0~���B�i�]�u�SS?~�sx�t��K�Nz)�0�C�7�_���Uc	�X>��[7c$�E
.��d�ҕ���竸 ���9C�8�����Q�Vrǜw� �0��.4_�<2�>iȨ�K���H��ޙ:�֋l�R�	<�`�f�%�Sh�d��"���t0<_�]����`����9�v���xE���z���^�ə���&�#Ϡ2OC�f�3����%,�*y���Yۂ��i'����kh��9l��������6 *-��3�n�׵���2��졍䮕P��8��'��@^+U9X�p�)r��&�����XPI�eK)��O��/ I[��#pRH��2]��r��Ȉ=�C���H�DR�Q��P����5�|d� ,���VI�J9O ��t�'&��V��$�:3�U��Y�G���)�S��N���T��:.���3l�S���y��E �n���<}��ė<$���!B��_a_�=6S�����B�QRC�=|������=�I��"�2�?�a_�^��Z�d��+���n��
�Y�T3'�����Wn����8�@��焚���c���zm/��N�#:Hf|��4��8�~����$q���N�e�+h��,�G�gH�����k�Ƙ�i(��� ��b"z�V�:����`E���*}�:c�%�|�O���q��Ə-�Ӵ y.�
��}�~��P�S������XD�
G�J}����>|rTKēÚ9��]�H�� �2[3*�1��1^�󂁨�h'�M�� ������mz&�flO���Bvd��:�nf)�����y͢�5���sI�y\
hɨ��]�O�q� �&Q��Kp��j���u���
3b�-��K̢_���r�Ք�M�t��K�ۈ�X�f/Ѵ� Y��4�� H7iE��*��[�%��&q���n��sSY?�"OaY�	`Rom�O�+d�o�H�T�)��=�K?��J�p��[^)��n�|S�1��,�Xz ��AU�6�k�FM�r�������Fۙ�5VM׶~�����2�S���n��{��f�8U�z4v�P���$Ͽ�6��������hG�h�K�YJƭ<�L����X�z�_A4�����sZ�b�L�ti��s�[�%L�c5�f?4��"�9���i?'����g�*��|�_y���b|�����Ý�WkK�����s|���$u<������Ju��hX�y�5�f0��k�`��|_��CVQj��X�H���OV<��Tn�s|�Y[� ����p/���=�Y�I����L���,]�N���1��`��1����ǿ��Vt�W$'(V䂎�!�[4�L��[��c�)I�_�o����4�e�S������@��*�����)C�mkH�&l�Nwςt	�]���dw��������G�[!��J�i>��;D���#�	#>��������"�;;��N�xOq9T��Sd��s�+�'�쬈񹯴H(Qb�Ϸ�
��ĒkZ�XW�����U&������L"���B�$�F��8�>��rn���8O}y"񑖑[�E�z���na��7}���[^>���zh��>�����9��JP�nk	�unu�b�i�����U桂`E R�Y�ǝ�n�D��8(ݩE)Y�u��֮��	�����׎�V�|�,Vl.WY���i?~^Rd�5� �J�^.1���k��b� �.?:f64��a�@�|k�0&N	��_<n���c����< D�=gɨfm��䣋�Ђ9�ǧ�u��A�vs�+ �(X'��g@z,�B��}�e2̯���:�u+���WJ�Tn��d��g�W\�d�d~Ҝ�7�|^u�e5�ؠ����ѯ�,|�u�}����WĖ�M~vl<�U�yK���t&?�A�3o'gQ��� �_�C�e��&hT���BM6�����F��JA��l`�yH�b��k�}��0���.��,Z��!Y�D�\��Qzc�X}��4Hڠ�_�}M7Tc����bѡ�=�hS��؆V�Y����#0�+4�����"|Q���("6�1��?=с:�9ƥ-5��VS�Jx�8�t���^�OZ��:�_B�a��|"�M��z{=�}�mD>�Xdn�9k��OU�`j�7����(�{ޗ*Oh,��x]/~r1k튞�|0,���J��_w�!�|@X+�������h�t���|�pGB1�N�sb XN�n.W�`�1`=��&�w?�e�!C�6�	rF���Nħ|Q_jL�Z���ڧ>��V"!���Y�9�ѷ���;�1�]�r�ѕG�*��Ό��=@q�c{b���R��>��TU�Y@��塃���Z�	�x< �}%&a�%���p���ԱH��&	��w�ȳa��XH�f����a*%��)�:*IQ�\v�����Ӝ�a)$�������3>�������� �/d���ə?!A��L{H/�b���Tw-��S7�	��۷����]D�끛ЭCb�Cy�����Y�ğ���@��ybm&�����q��,�U�^5F`Mbv�il�Ө3P/�/��j�g��_��ο8)!"��_����r��|��>zM�?3�E5��L��Ɯ,J�f�xo���Z�?Fb���DQx�^:_>B���'�6A�0a��Yt손[B�s�r��'|]D��alJ�D<��,�u��<�ʵ�(�GUc��t��L1}�(q:��-�x��7�,e�����^�����'��QSB�ѱ|	#]V���E�	>�iy��pb|In�˒NU9<6�	Q�����9.���M`yJ_�{�=�#�-1�mu�5}29�t�a0X؝��M��̙iw��y���0�!�a��-�c��7�C�"�>	"f׍�p�s�|���Hn�̄us���vi�hڕ����_�Pi�5qw���Q�,)E���0���o�a���>)d�v2��2Z���>`.i*�y�a���Q���h�ky:������B�΢D\T�T�h2q�l�rH�{:kmT�!�9Gt^�.1#���6֍C�n30����Y�!zһ��ch$��7��\��߷x|��9L��D�NGl���qo�Si^�Ve�t����ƧA6'4n=�͊[t�S=s2ė�%_�G�>��-����9z��[ ��n}���Ò�̸q�� �2v��غǅ�Ѵ��P�?�A��a���x�L��i���k������xƙ�E^��Eç���VK���-i'���c�X`/��ƥ�h`����8���9��z(��)r�}�N�&Uϧ(�ӵ�=���FU1�@�B����"UTې>�;Mǧ���r2J�Q/�~�{�c�Z��%
	�4/��2@�Pϓ$��)F�1<p�<i� \���)���2B ���D�jB ��'����˫�ގjոB��/�S
;�E����G�R8�c����RRS� 5c�d��4��q�:-�͹Rr��8�-u��Ĝ};2�;�7�|V_i)��eY�X򤵦l��\��l8d;����ˎh&P���ۊ��9����Ȼ	W&�MT�CD���7/T��\�=}����=�E�3��l~����h	l��ϣ�`�@�[����� {�.W�5�/��h�)�h��=$����]"Z[�ޭ�W�vl{:��n���3{������_�B�)�������3{!Ȥ�O#7Qr�2�ݭ$��S��Lm���ښ�ܨr�ڿ�
'���#gޣ�4�X�*���Y&�@���ҿd;����I�� O+�&�r�y�G���O��
;��3��vW��B�}1g���nƷ;�o[ç}��ƻJj�C��B�+�6٠���`ؚN Mϱ��C��02��.�L��)H{�oQ���X�Ͷ�3�G�J݂��-�-���7���뤟��Q�����z�}�ݻ+/h�`F�v��s�g�����-��_��e]-R�2ln�(�=h5��Ѡ{��@��yB�������X'��qtW+��1�~� �T���5���тzƤ�Z�2"x
�k���6)8�0���2?;��Z�G�����;���U�$K$���!�c������]:d���Nr�LH�*\�H����.A|Q�|x�0����O�{���sU���|�z��A�N�4G���/!�� J��V���%O�z�(�п߶���p>MT93��:�f�:���(wjWF�9���D�Koi����K.�_�U���o,���$�)r
 ��z?��Lo	Pll�(��?O�\�\3��~vn�.�f�2]V� ���.����i@���L{��u�F�����D��9fý���Zz+�21��t�V�c,�����q�D�i�3����w��>b�2p������!q���>��O��������W������A��~�\W:�B�I�L/r��P2�%�:" G��*>I	��J�F��>��I�O�|��_����)=�F��@���A�G����
�y�2'��C	��	�(��㟸>�?��--x�������4_z�
�`��W�R����o>���i��}���T����@��Hh�B�9��8�Q=RjV4:~;i�*Y�b�G�ֽ���(���J�)�܎��k]��$/�� q�'팚�Ѱ��G<\����nO܈>?�V��$� Rv��8��~��W��
�]6haR��rQC��M�,Ju��O��>N���C����m"}�S�R�J���w����:׽�$@#����+�^Fz�^�P�0pF���<����\F�;άge�����}�t�s��]fnYw�9
�٪)���mLq�g��q|�V$�Wu/n xS'wR�=׎O����}E�X�Q /������7	O���&��)��e��ʃ�CN%��f��!��ù�a�ց�L��6���挘)@H'��m؜4�% �.x����u�iְ]��Y���Onx���|�@�ƹ��Ӫ����^<���u��ͥ�*�>�eI�E8f��L@��,��e&o��B�3��k|���C�GǓ�.	�������o�z7������R Z�[	����w��4�ކ%�N��Ȟ��������H�,�)��Z���UM'$Ǆ����!��N�n�{WI*ݎ7�E�`���R��N˴���m͂I� �U�?�	13�N����ɐE|_�j��/�M���d�N�r�
����U����1Jb�:�\(�q�fg''�7U�����լ�:7_UW���f\� ���{��H��8��/���D����G�U���fO����)��%��v��\���Kf��?@G慐�X�&��!�G�f�*y�-ئNA��Q*8�����e_;�:�2Ճ�2⋘�b{u���R	�׿��O�sl�G�Y�ZV���Њ[�t��A��Ȧ���%eC(A��[�GP�<�1p���p7����1Ԛ378mN��蠻E�=�zP�>6s6j:J�o@��G3UM����n�.Oz	�1+��y�+Ղz�
a	�m�Km�6�e���D��s�5�m�ge@qG;��[l�����I�1W�yL�=}��,��p���S�D��t�w�Ӛ�HG�R�ն�O&���h��]<	�V��Ѫ"��·��=&8J�0ל%�����D�Q�c����`7��9c�r��ʸ �,�,�P�RG��m7�*����{8܄�%�tO����k��VIVD��(I�T�[�;gb�͵M?�mb��e��ᦏK_a^2>���\X *�89�����\���o��oGfp��bLp�QU���?�.�@��
�K2}6�hK��b���7�N�C��0�5�4Φ�o��5�r���Mg��a��3�"�0���#��v"0s~rg�����üAEX1aPi��R�O��@�P,F��Ձ뻦{S4��޵ vTL����,F���$Q�wx�����P���k5>:}��NQN��XYߏ���D�*E������8	��$|�m��R݋��o�7�,�k/�Q���F։)`���9[fRp
�&�����{-����R�M�_��u��}��ϲ��]*&�����2Yĥ�h�c:d��룒���
�s�:�vc��.`N��J�����z��j�B���i-|�~R��|ڦ�Uf�E�Dx�QB��>�IH�t���,�S>�$�SԼw�4MF<�&C�w"4��v����b?N�c����� nK|�HCq�g��R~��Ȋ��ʺP�c��u�R��c�'�	�8�V�Y�6�������(�kd +�p�p��[/)G�����7�kl�����zu�T�J(f�3�q����c������e��)uDI�^v�T�]%7�������#����eCc���=��I�1e�htFÄ����T9�mX/+9���G�/ዠ�u�	�*R�(��(s3�����Ԝn(?��	9��w;�ǲ7��m�%�hH�'tk��~��.�"}X�'�cc
���1�e�=S*�f�����.T��=�4AZ���w��5�v�r�{�Jz��5~��/R���]~æ.@
{���O���,uo��k��w%Iԥ��l�O���5�����SF�X�)J�9NV��C�!���?Lea��~aGkE~P�{9h��*c�!Kc��es��=���^�h5.�$���^���ݢ��K�/i)3ٗ�]&����K�����<풻I����`8�΋�� , �nx�Mxѹ�9'��X�H���s'�o�7�E� L`F�=��NS�Pq�� �c�;�����֓�;�3׸�)�e�rSG��K�+B�rUL��_A�X!�����S5@H������5iJ}U�b�k�DDH� �e�F���w5H�<mJ��^�}M����� ���Qxc�(��=�x�R6��N7�^�(�rV\��"	 �f'v�`_e�(DDxL�T�}>��@BL�J[�P�ף�S�50�僓;GC�颩��&����~��M��,��5ӎꗽk�$k���$�./V��]c����5�[����s�m�[�9�h*}�ZM����TR1�#z?�R��
�3_��:��V�R�Ot�Sct��Z�	^���,.��,�|�G��$����w}U{��zA�o���;Q2L�&(� п��>t�*��w�qϱ�5�z����mJ�i %�����z_ �)%t�sV%Ʊ{^#XʁÆ����R_zu�~�����/��hV�6���2���`�h���f��5ql�{agF������4:��/��[آ���߶��\�2B3?�����<��$�wΚ3�g�}���[���~Z�S=©�X��q�I�6��^+�����ޗ�L*�((О�z�dUrHH�"���e. �U��筊N9Tl�q�������	L7��T��p�'�mrY�D�[:�_m&q�����" �q�Dî��x�W�'5���
��[G�w��UW7:P�S��4E�[]_V�|��	��%M�%�	��r�o�,��ؙNs	��f��0�׀C'�.(<}y��b�o�5�,�:�4��$JJ�j��m(X	cjd�u!	�Z�v�:^�P� sԆ���n�C�!i�{R�K���yp{��b@����`��I.9.�sL���]��ᶐ������QEJ��#��:Z�"���R*�U�M3#_��"T���M��3���92������bz�.#�W;G�)K-��-��%f�U������8:v�i.�D�
��myiSUC&@l̥T��@$l�1�����(����x&.�@%�{ޠBMf���)�R�~�M�]�0ѿ���w�}�h��Zcd����t1C���$�44ܺ�wR_�{�<����%�t��b��� b~B\v�~�c��9���ㅕ���k�
��3�����\�UR5u��0vk7}�}�#�+�/i�� ��x��h�n�[n�}V9���A��^٬�23-�(p�&3����Z*��x)�����h�}%��G�Az};���!��:_e�@%���~z�����qm�~��KT���E��/�)�Iԁ�.�;�*yi��1�3��TH���{w,���c �1j7���H�͏[K��v�Ó!µ]bQ����ԼW6��1����uM(6�"N����u�(U8P��<<���0K��+YQ$�ë��i���ǧs��ӱ���,�#,��Q�C����Ej���#�z�F�I�����p:6�K��68�gD'-��[�gU,�f*���AK�MI\�R<���� Q6���uK�Q"A5�v�<��O[�ty_7�灥
<��{G�k)e�/7�2��iyF����]��r�Ysa��5+�R�34�{EEc�j-XB�٥L'�ߗ��C���Uݢ"���8#�����t �PYKBۂKO(Op���2J����{�܎}�����Nã����*s��*�%X�O]MN2�`��R�ى���~K�%Z��,�Ъ����)�7���B�y\{��l�Yt,�*i��s?*d��pͼP���X 5� ���8J{�~&X}S�-���CyOF>M���<���-�mx��X[*GۈT+�|Ԉ0��}Y��>&�.�N�����?���h5*6��m�9��b�y+%����b)J3�^��"H�7J��S zvdѠ��y,����3�j�7�f_|��M�w銩��SK;M�K/h�|k�b`>aQ�fe�d.>�@���-�h6�~�g?�2�m����0�ťn �(BN�ay�o<ʺ��17�%��o|�����#��"��k������3}�A���*�udi��厯����D- �ۑ��m�������&b�Q�~�]������ɷ���RĄs��X��T��"��?e]'8!<�p
Q�W���G�7C�k>bT�ML���R�a����h�"GDA �w��`;. =op��	6v�<˝�P�ǎ���P����w/W�N�8`�#�D�տ@*�IZ�7z�3��\KW��ݮ�Ԏ�A+<p-D���&�͊�ӹ��M-�8�Y�
�l���G�;��n��"�ݻ���m5��I���-e<V9��{C�8uՎ�Ltx	��;E��?��fµV�a���ם�~XR!u�����37��(��z�ώ���L�,j#�J(h��y��l�<[��/�&AS��{9m%���w��8b�(���[	��a�����`o\���,�Cl�&�+�Jr=d%�����'l|7B�;��ISՄ���wc
*��4�~��PȬ�	����l�#�DO�gv���JЄ���_���9�Z�p��Yļ.d;�.p�J��F&���d�	��%ZT�Yq��o5R�l�2���o6�Ϸ���T�Ƒ�?`_ԧ,c=��Z$!�IX6W/�����=;Sf��2�2#��S9݄A��%M!y��U��7����hu#�>2~�K%zf���
P�&��A��h�[S��}��û��<�����y���XCA~���q C��p ��h�`ңؗ�����l��hqFUqgFd}(��^�ޑh���^���A�g�qn�h�����6Ǎ$�F���(��~cAק�ʲ��=�LE��S��!e��H��`��Ǵlˎ�R	H�d}PX���Ȍjӵr�%��8d��r����t̩ݺ���1�*�z�췰��b��)4�	��F���׃cƀ#tF�p�bS�s+�e@7�wX!;m�ї<���s�����s���ew�@ۿ��_#�R�)[���&��]N��Sv��yt�U�F��T�+�����L���j\{�Jd�ڠ�3���\!����C���C����=���	�.�B��Sn>@��W<��d���1����VBm�Tx� Y���k?�4�wv݉B�-Р���:�4t�oZ��d���l^���ٷ�����KdKzM�_z��X�����$�v"���u�xK1yt�5��?u�-�9�=��!a�MǞ��f�$����25S�/k��Ș���0�/-2yu�zj�}�ß�n�G	����q÷�M�,2>

��>���U��A
��V@T7���p6�Fb��S�uW8 ����@���^ ��3�0v�i���ͳ��\�)�Ef���E|�?{�����녂y�;����eH."��Wy<��G'D��
e����:
9au�s�5!4 ш�K�.�}0a���� Hw$��[�L�Æ��3jx	�B1�uF���d�b�?��-��\,M~�����7���ɍ�4�%��XNt�&�f��O�AH�^�Z�t6�G��s���gI
=)M�$�ј���`�j�����8��(�`���W��H��%M��n�
h� ��b�H*���d)G���5�������\g͆c�\=o,G�d}���$G��$�ge�tJ	ޠ����26�	5����m!��i�~�N��W�p�i��V,��;Kβ:1x-����F�O���</���C��d���M-�
�,׉M���M��k�X d�b���y�q�fb�v�:a [d�v)�05U��=��F�v+�X�
$���=�|q��Mȣ�ŕv�A\��iD�3?����C�d������a�N ����JP<l!�����|W��]0�Ȕ�֣���a��{��e��#�S��~1�~�F��I��RG���$���w�zS{) �O��X]0���nV���ug8˜�%�in�^��qؖ崉��FK�����m8�KQR�J-�N��o����h�T�M����|���%��iq.�-�6�p�½��۱�R��W�ƷE��c��0<��
h���$�T��0�k�P�L���H\��cU��Qx�k]ܮ�*�<�A �R������m�����3���o"Z�Dc�� w'o�]�3	��o������1��ްZ�gU�Lv��Ϡ㩝���K ꆛSj<��oF�V:��T�RD�s������'JS@(W�-+'�& }w4���B��?Knp���S�DF ������S�+Iľ8t��ѥ�_|Env��@&��܌�s��R��ߗ�4Y�п�f��.���D��j�gy ��A��1`�a�F�|��Ng��`l���4�b}h{K�,Čs3s8�z����]���*�k��ޚ�<��o���^�i_�׋����K�K�x��I3G<f��jHt�?34ߕLv�2D��Ԇ�;�z���z��T?p2�$�."��i��G ��D�@�8	�@�I���T9���!r�ֱt��t)�=�u��\�Ös:W{NtĪ�_���&��u���ҩ��2�y�4J���:jf?Ͽ���d|.���r��+�k!����O_�ѯ9U�M$r^��I�-��mJ��]��$8?T�uh����=���t�FE�.£��o)�вD�;F�^1�l[����#Y�YzI��ivl���@-/gn������T�FT �=עǔ�m��~���9�_���68�r���b�{�6/!����K~*�p� �����ղ�Ms��hXx>�a�f3{��`�)Xm��j=�C�@�
{�D�V���/e�x�ʧq)�輓״˟0I��]e��]ʃ4#6��	?�ByP����:��獴�Wn{",1�:C�Zs�֩X�2$���3�6�&b��`p�@�\8��'!
؞���i�B��ȱ�Y�6�����}_���"�v΃����� ڥ<-0�(���1�X�U��U�~=�L<��O�l�5�f(Ct����ķĩ`�9֏����'3�r_�F� �(B�S&��_6��n���e������d�Ȕh���?�
��~?_�D�D�0�y���ST�N.b՚=mE��+�%�b���q��Q���)�ȼ�X�UY�m
�[7��=Ǹ�'4;&?9�q�i�����㣾�L�m)��I:����nǊ/6_��q��� ���[��j,��9~��rfq����g�����O=�
�>�6 	�����Y��>1�H%�"���ΰ<�A�wV`�m$��j1p�fm�;�T[ƽ���1B�^�%�c
��lVJ���b������E��!�)�)Qr�R����iƿ�	k�!�����z�����gJ�	����9sy-�h�T�9�7�vo�Y;C���=2���׋%�MjO������a� �Z��e���3l_y��H0�#r�ۉ��뤋xAi'
�+B�*3$23��Pd�hOU�X��E���M<��Xʈ+�-�ܹ��8�|���L��ɡ"�qa�y�%~��YUtϜ,QUe�� ����w�T�8�&���?�8bӝ���zr��ls+y$�[/x����+|��Zl녏�g��O%�{z�ܫ��#pevy�-͈�y؏@�*;R���c�b�2L���췘t9��#�H�?�Z>z31L]\*S�l�!���Ԅ���
���=������'����G?'�I��Y�<��3|�|�;��PKA-�83��ݭ��l,w�9�A�M���$���,^���?��_�nf!��(��^R�BM�؅J���>�c�[ ���M�r��Ӕ���r�6C����y�+߁�W�"�a>o��@!���!�*s_�?�L~�0���l�~磒ˠd���=ԡ%'bE'O�b�=Y޿�>:��t���ˮ3�� .F�W~B����g3�/z�z�6��ȣ��9rJ�^i��U�x#�73�`�F����/W՗�~��6��j�3WY����jK�\ o�?���9�X����c���ܗڨ�8Xt�g3!�J�,b���+~,iuH��M^g[Fcq�/Q�!z[�~h�aq h����]�����ޑ��|k�9Rm�̨0e���|+����2[�{I�^	���M�Y�Y�n�Ա̄�d��u[B^`q�V�|�齩s��#Sc�ɖ���9-#A���fX�y��:�� ظ�'��0�\ؿ5����8��_��i�D7�KM�(yy3ɇ��N�q��R��>e�Q�fς����vk�9ȩ�O����l�ڶ9�}��ڢA��a�J�(�@19��
���+<@1���7Y1<���1�6l�6�O@�W��<�h�m��<Ja�[
���'Vw�5���W��4�!.�&�K����e�M�w]��K��p��:��[��bIe�f�>��	�@��ٻ����n� O���NSd��zԖ�f��]�0�[bJ�qֶA3S\QC�Uq�m�5�6櫕~���P.�?������b�c��?�7φ��f�"�\�G�P^����zmg*�����I��R�7^�&�ㅈTF�(]d��ߨ	)�|L�I�D�A0��r�0�#�M4&���h�?U��j����	�G��S�?����Sc��<sW����K{A��e"�D�1;_yX+�V��
�LBV�%���}��(�愽JT��pa��Fy���ҁ�D����n�������7��$j$��#���D6�Y�'��o�r��ʓL$��a���޻�_�h�z����i!�:�Ns")��ucS�~�v�ۺk-�*��(y_����-�d�!ɀ'd�X~A�n��ݓ�jI��f�N9&0re���$��	�ű:���Ě��]^��_�`62��vS*���s��o�;M��$1��K�Ճ1�͌�n��� �y�@<�=�%�qKH�B5!F��i^@G�3�S/�8��1|ɘ/�$x\>����q��q��l���|;9����V�|�pY_���wx��ʤ�B;#�������#�����p�LF>��G�p��Ψyn�bJT�H쌻�G�g����r� c���V�&ZI8�t�� v����L��c��� D@e`�K��U��`nTAQ�؋+����av5��6�hl~�euB�0�+|�"!���E�0&~#̦���7�ܖ��~�p:��\��)�.��Z_8��ه$�l��!�Ef)J_K�&#r����8�V�:��]>h�fnI|��^�.�x�pNϹ&� d޹�����x|⮆���q�c�)�?��3@�fJp٤�:U�W�N&��OK5GN�ś=٘⽃�I4�b���-�8�U.�(_�;_{A.�~��Yj,ֶ��:s��1�O�
���6U�ۮs+KUM���ע�=�0�IӤ���_��;�eFy��@�)=&��[!ZV:��0Лa�s4d�1� {�`�>b��@S���-��62q�o�0qr/�b�[˝����?O�']]JMmpB4��	H�,���fi.#�k�U�o*��Uj����N`��2���'���_|�m�y�mէ��S���Vz_���M3�+���(7��A�[�2�Ba�$����l��9[>q�1'�"�K�|�O���I2S�z��==��ǳ�m�g
�cy/�!>^��x���6�Xx����k�^:���vȚ�|�9I��i�i
���k��b�H(��^�㜁��'�L�`��?T���c3� OP��9��k��n�9�'���12�~���U�*�R�ݢ+�HV"X~=ɝ�t?Vb�A���l� `��4�~��}�*�������pD�0$Gj�Ŭm��zQB{}��)�b��e�v�V+�Ɨ��8��B�VH�uC���j�?���X�%F�Dz7����䃱TDw혀��l�%���<�����}E"p���.^RA�T�K�D�!F�gDH��,Y S5��\�	0��@�8B.+-�G$�ȏ�ya��QqYR�����Z�I��m�n��Sӱz`��v��>R#`��:�V�gI���'��bb
�@Kҭp�|����op���k
��¦�����O��>���R��
;��+�[��IP7/|.��7�z"]ՙ�^��-��'�[���-���/y.�P>w>��@ac��:�;����;=��&O]��k�� 7���a�B�
z��W�U0�2�h���8(�eE1+�{��b���dJ@uk��� yE��r�t�5n���4Z*9N^�P'��h}Q,�GZr�*����J�2����o �+���v^�GA@`��?��<���Vu?Pl�	��dc�-�!-a��U�1��$��)
�W�_��;��^�O�}�'�;��
��q�ᢙ��u��t<��Fsd��&��eH:�J�� ��N��]S7;��Q����;)Ue��d� e0�@p�YT�R�k����a9���ޛb��RSPg�����k���C~����[��2�Rk��`�[J���9�0�#�����S����5�^J���>��+mȧ�UxֹZ�6T��|@q�A�LX��O�I%Y��-��_38�����P����M���!�H>��i^衑��I#���B���cV���1B]�C���Cd�\.^�_�L�7�b���Y��B�"��p�r�OZN���[�V��*��Sܐ��,�5z��è��0�_]�ǒ���3�F��e[��6���!���0��R��ya���E���w���#�l��9]D�O܃.o$�gS����9l `!��tٽ�fMA��$�%^�����(i�*�:d���V%�u��3t���y�~��V�e�js���#ȅ^�6�jp���83�*�g�$�o/
���N��$��:t �p���v0�$c;�1U�9�h�h�o�}8dj��
�լ��X�'�
���� �I{W�>O\�Ʊ)쉿\�iH���MZ��ë!�d;�^])2��]I��h�6|_�E��^�]3�a����Km��(�w��*IPf�X�j�E]-�:O��My�JePU�O� q��%�[�K�o��U��g��KJ+yHܶ7��*��㤞lx�b� X�؍�y�a����j��U�ݚ��b�]��}��ؗ��v2����0�	�P��M7��U��'-��)[$\mX�x�/��􃳤{$s���TR���}Q�wqv�m{�׃B)н"����w�Թ�x/��Ɓ�W[:T���S-|_KFD���2�� x�,{>Φ��u�xb�;���9\����i��r��3ŇYl��}�C����<6�U�1FŽ���p�ZzMLf����?s�L�,��g[��L�ވ����9=�m��q�)�Y8�x +��'\/�%>����y��O���!�@��}̄�늣09�NK��⼑��~"N���g��t��|yX(`���KPE�Z/��q*L���,����1���L����RZ#mfȈߏ�<D��F4-�Ѕ���8o�@B�Mva�^��G���|��䀍F,%��jiᆭ`���Y[$�-��A�����D"9ҡ�l�00�/=�y�U�~���'S�>oZԯ}����2�RZ5[޵7�-�HmˇqƊ��O�sv*�vͩ�zl��҃��rf��F�OE-��*�8�PƖ������s�Cp����;�bb=�O6X�������5����D���V{�dq�F��'Q��Ҷo�é��ղb�p%�T��VbʷY#51�(��[��SM�vsLkԦԮH�o�E陜��X��qQ{�0��v/��V�WҰ�)������.�ҁ��|��a+qE��V�6�	t��F�\�{� WC@"��>������ |��S/ӫ�<�þ��|��?a��C���nײ�Bߒ`ʝ�� ����8ȼ�0C��*����N{�4�>ȳ��Q��g�PxI���(J�Y��w%|��^�)�g�)͉�!D"�1}x)y�;?Z��n{oN�I%�2Z>�&f�T�B'�ȊFʹ�8ސ��M��%��
�i'�C������������5��(��J�V5���X��aj��~c�4��f�+U����z��
���������M�梊T4����do)���w���?l0��۞]93��������"��U��|.�"�wX
?������q��u 	J��L�Zͮ���$�Uh�?��X����#�2&�ߔt�����d�����\0ݕ7SDWI#�~X�$���W��]�!3�Xt���RO�Ѭ�8����x� ��J�'��b�CY�b֪���W��)V&�RM 1�c��%���n��O�{��� �Y��!n�M#����K�r���FMټC�M�0��I�C��٢�1�S�|T��o컩�^���P2�{�J���CJ�WY�B�2���+�E��y��x�pvA=��F�<�a+?�V�d~`I�{l:O��N����_�;+����Y��N܄�ra�2L�3e����s5�ta�,����-���R/Մ%,6�����c��o�6�-�_��Ǵ�� l���t�I.PՄ�����Y�`~pTzH0��u�;{��$��O21H:���Z����`��������z���\1���,�r^A��Lś�$�zDP���..+<Ȥ{I^XQE�R�8�ʛ�c[�
��g5����%�������zZ�F�`��	#o����U7��a>/
�T᱖D7+h�7u�SB�T@��zʓ�_�+�$$��-es�q".	����&N���m��L�H)	�Y��r��9���
����2��t��C#�@@�����m)W���	#��s���F����LHV��nD��ٌF��J;�㤈:'~��F)8��燮 �u�y`���7�0��,v�h������mT�^IF����������|��d��r��I�`c�Y��Z+� �(�?J0�UPg%۹֑]�v㇯�${Ő��=����*V��2��cG6/HjZp֏�j�X�/�U�q��5�=�ޭ@q�J��c�]e")��4�G[ n^!x/���xoN�@��8�7V�b�җ���0�VE+�;?6o�3��6��3�Fܣ���ɏ�4ض:	5�s����u|�$�<Rѱ.�	>��	��%�x�R�8o��˺X�!��!.<Dn���	|�sF�F���y���b�8���AO�������`���Q'�QK�&t?��^D�&uqR��\,��{nh�@�����]��6#�"�V	#��!��
ڟN�;�KYdTN[Hir�S3���8�ʶ��ԲH�����,ڎ�V�8adh���[���I)B|5�i@�0|�Ok��X@d:����&�E��<g�>F�C8�g;��ś�<�Z�_��
���8����ݥD�,s��#�`x���.m��\n������5�9�y��bq�U��q�@����hy�x\c�`��iK�����m��S|u�{3G^��*�&\���ڕ���+>��݀�p�SGʿ����^Hq�|W�����=��<y��[O�?���<� 2<�Z��u�ݥ���/u$[���C��K��}����9o��`�*��%J���������a��Lm�)�8�5�;�MO��Ƈ ���C���Yw�i}9�� p�gͧ_'�f���|�Z(n#��dP�gε���+���]Fi�M���A��T�ѧ�OG�#�e�����eCmRP��E�(	�FNo���x������Q���N�h�g�%�)>%�>�v��~��5t!���Pe�*(���k��F�F�'�$&V������&�C��� �������T=���9��]������A(��Jg��%s�� ��l������4An�J0�Z���M�;=q���o�=\��wq�&O�"}��������"Ѷ���r)2�9 �ܡ���ao+��\��U���#I����gG��џ�B�m6��4]Q9|���K����י�h�wס�J�O�� kr���G��g�n���b��X'������բ�!�Ά��X��i*�v��Y�7���,dG#�Չg%��w��)RK_v�*B���zp`eTut���>G�/	���:�[$\����
C4�Ca�+:��4R��cj>��1a�e{�ۆ�dN��M]Ɏv�$��/4+<,͍ء��(��08bHyf`t��^����B�,���"�%u��ho9��G�M�L:������߁�)�B������뒾�~���f{�b��Q���NY Z.�v��8�w�֗sʞ�>+�i�b��J�`~���P�l/�Լ�i-���54��n��5uٓR	��i?�S����q�H����Ũ�e���ޤL&�E��{?����L�ҋ.]��\&ifS�F���K���i�O^��;��-���NH���N��y���P�dB;Љ��@�ZRe@�Hq�j��_>��З����]�k�� G�gҿ���Ӑ^���3C̕�|'/	r�NIJ��`���:�D�/`�c�yly�WU|~4����j���w´8�C���/�f��B�꧴}��_��.΅ɼ�7Gi�I��8��7����V_����(��_���nly�P�WC(�q����X^M�x���N=���f���
�޼��|K���V��%�Ǧ@�̗@q��d��m�bB��}l�����{��H�v���N�]˧ο���\6I�����e}h�Ŋ=�r�)YpS7��+Ĝ2>���p���CX�����&�����؈��⬂A���)��(M��ݦp}��Aڗڡ��1�~:>��ʑ~<�֑�a<Ϊ�W�u�N��Q=T$�5e�$��ď"��e?|�fs%7��Z��B�H���l�=ڵⰦI� R�{���M�����Kؠ�|3�r�*0G1��D����.1{��m��l�������4��+=\߲����l N�{6��w���d�?"Mn�=�Xw�9H���T5T&�]��Pb��\'~hb������&�R+ڀ5���g����0y!ĜS:��k��x�j�u[��:W��Z)H��ڿ갺Q��y?M�]�V�{
XU)��g���@蜬�P��#�۟5NǪ�܏���I�l >��#zl3q����.��M�B�xwj?�QFkp]���[/��b��w4�雾Q�/q�w�:K��Z�L!��Ռ��ޘ����y���+�t똁N%2�YͣqBs/�ii�5��1���e�Qb�&)�#��+2�v1�L�}�ͰD�4 sي-��A۽9�K_��_.ږ�f�3�^;�g������dnG4;�`	�{��THd���4f�"&��(>�4|�ૄ���e%յ���)���{�xMQ�d#֓ɺ�\�c���s�>~��%[��#�@�7�wp�6�,�Օ�ڔ> 9gr*	j�C�=��K6�~��z��Ľ�v܎B�&}��.���\����׍*�|��v1�Ȓ�E�tޓt)�Z�B\B�u\ #m�k�Л	�)��I�y�3\���V�X��V[����3���y�hu��/h����ZO�,��\�M���mT�P�-�<-���~<�\��!.p.� +t��y�e�spǍ�e��p�o��Aȼc��vƐ���w�$�c��P�����/.5Jx1�R��y_r}iq,�b�E}��c�+�Q�nAu�����=jWnE���P_��y=���p���ZV�\��)�=x��J�z52IZ���j�q�B���u�u�̉^�5�!�=��4�%�D[��8�pUՄ�t����tM��(%���~��E0�����W� Kq�qB֎ky�5�Q"֦��97�����w�j��x`ޠ�~3C�2 Kt����z�!���N@�4�1��+�4W]l�<�k!�~�msxn/���^z������G�` 8��
>�t��P�i����̂�/6M�U�����D����QcX���e�{ɦ"�L�*��P�-TB�V��Ơ��#s0���NjN5�T[Ne��GېD$X�j%�3|��X57Kz��� 9�	��ݟ0��
�_��)�Y�&*O#/3U��H���	9r+0���ܼ�~�;��@n�8p�e�D�"u�{���}����z�;�Ѱ����*o��(�~C�4�|⥼��N���d�8Iv�b+_V��T1.�����}x1^y�d۠ `�L-��\����)�;��}׳*�#�&;�N������T�{x$�~�a]�8�Y=#�I��M���YI �#�Fu�Uidekiw��ߥF��`MI�?(��(�G���z�_k͢8�gDuR�9Mџ[ظ��f-�����/�zzg#a: Mt)viD9��Ξn�ӢO�9���S�<ٮl�Q@q��SQ3Nk��,�&��?ps�W�0����]1�u�e����_�3iR�=ͶbU�۫��Y �E'��N��~*pL��z�)'�া�f��7܉�wq�?��@ȍ)+.y�.��8�Q�mW�K���t��'��%�"�G�������LkHN˾����Vq���B}�&z:֏O@�hul��j���Dhz����MV��/�w�>��ȇ8�-+qB��KM� m��@{V�땛+��{	
��]�<v��r�K�_]�z��7���(�2�^k[
���υ2���n�ͺ�~�7�X�ˉ����Wy|���Rf.�tS}�Uh���ڵ�V���en)O�����Xu_��S�����������]�vst�d�xrI7�O��F/�ǣ&]�<Ȩ�lv�"|6~)'U[�AB�=(=@�S}�+��O�փU׸x�kv�f��c 䦟z}�g�!�T@nf
ݵhV��Q��2��2B��fx�]�Vz������������B׸1��p>e;8i�1��xqĞ�<S^/{�l��d�m�<�\���׋�����"�kTÿ������6��� �t$%qV�)�Y�EP���	(P.��t/g����J��n� '�ź��<�F�)dy���ģ�Vt���*���=/�\t���Y@����%��Gi�_�y�y���.Vs?�֮i� gW��-S?a�z���i����V�[6/�����V�U��l�(?.H�^ږTrͧI�5V&5���� ?DG�&��Lų;�?�� �x�&G���"�pdv��.�~�p��V������m��w�m���ߐd�.d껸�<�� � �*�e���k����a��˿߮���Q���sS��f���C�Ʉvi��4��!d�P�h|c�k�RկA��Z!������~Wp�?M�����b~햳h���T-`�h`��%�\W(h����SP4���CggzcN#U!M�_��/a���v����O�"hO�ԛ��9&��DRw�g�D�y$fil���X���^������	�Gr��_��{�e���a��i.A��x��'^2�Cq��[�!j�֠5�i�dŘ$�/84��5mg�]k6z�CT�����R��g�X7�{.?D^M>�F�M�50'�Рy&kITļؑݧ]?�:WL����
����V�ʈF��B%4���`*�V��JwM�gyi���Rs�?]O�rLy��;�.DNЎB����l��8ͷ�o�5�M�6[B�������4�Cg;o�!T�7�νE+1$uB'� F	�v��G�j�c.JJ��zB�4�,�IÍ��4�Nz�
\���?}B���\��OA?�E7j+���O�������<B ���4��ݠ�*I�.bpv:6�u�#�pЍ����:%���1��x��2\]�T|�"S�\BI���J��\�}A9$��I/c8�-�������7�
̀�GKTvݖ�|S�����q�?�),ZU9���J��m6f�說=A4D�n�|jl(��)O����u�Y�"%���}��P��Ĺ:Y3��wan�B�|<7="w��H���J�I)iN�b[#� N��J:�<�2�����S�6<R�(QS6E��N����*yLG���n��>tY+�"�YU\M�*r̍!��}'�𪧂#W��M�^�AXox�=W��n�!��x�U�$���>�.��Mk�?Y���
,-I5��Kgꗏ���!�0��/�jۥ�d{�y�`w�霬���G���Qa�e���H���5!&C��4J33G�b�����~�!�-��/�,D>��~�zH�;	���L�Yz�a����ʠg?I"E� r�Rd�|���吡)�u_f�DEo�T�O�獕�H �4�H%��Gκ����Yia���2&��o��$~�d˰$���#��,�R-M�s�TK�_����rH��ݑ��Ҥk�h�ڣߒ�T���༯�o�^�;A�B�,$������Y�5�������m*�J�E��Z����e���\"!�y��wS�����N���?ֱ.�I�����G��/@�Y_��j�%H�Ǵ�b���@qT7��uV�����^���2������84[����~�x�-��������#2SŶE�L�s,�<�<p87jv�_,�e�Ѐi�0�W:G�J�W��E�^c�<5j:��%�������<i�νLݝݥs��0q���{_�|�*���6�	�)dK~&�'�ek�"����G��K��$$$r�]��4܂��3n��T�͟| K����_W�E�����·m=NI�t��l��<UQ��w��m5�DX�����{z��E�<��=B��~�vu� �_�pV|�⑒�R{��W�GL�;�����d"YHт�w��|����aE��:xo��鍠P��L�1A�O����	��[���|p:u�dQn��B��Ӝ	9��ocTH6�ſ�3/�ug29�&q�Spp:-v�T�Cb���� �	�e Z�S��mw�&.�e�e�ʽ����I*>��s�����;ȸyfB?�����0�Nr�V0X�O���`��j.��a6����_�2ԧ�e\���d����o�!�����.�5y��g�m'���sڶW  �z��.��t�⭌��G϶�.c�(�I���/\�j�rj���A�� ��Ð�{����1Q�o�*~�@}^�ѳ�����[��.mݏ�=ͅ��|$gF�T�Z[�BK?��57nzg�
x�� �Q���(l�c$A��T�7L2l��}c�l��<D�Ti@�cޏ'���_�2"���9-=F] #�w��^(��m�Ѩʊ7{��߁�;��4aM
��� �l�����'LSRrn�#�32�L��2�uD=1�y�WL���,V13~�z&rG���U-�@;�J"O{��cY[\X"'���j�^��P�e�	�.����*&��6ݸ�ʴS6;j=b	'�#r�U��j�+Lz�UM���039��5�cf�~se��<aU�M�|��4×���n;t�L�a!E:�qD��J^��;�n��LBȕ�,'KM)mn���q?�,%nD�V��b�Sҥ�Q/"��bY�gr�yW|�aI|IXXWrT�)��	��+���G<�����l�4�l��EfQ�(����8�G��	'�;w��]EC����2�!��>��.���Mp2 �h�d,��=c���usze2��JQ%�<B ��O峍�-����^��{Ꝭ]���Ia��9vBB�Ɍ�˖�����_d��4��'��q4���	�V����)� ��
uqJ��\D�h�����;�yg��%B�"�u������Zz�V��J.�3�ޘ���E��w���G�:�&�K��5�U���Pd���҂-y��#�<[���޸�hF>��DX&�V Q��b�zY^\ըSr`m�0ؽhw�D��w���N-U������A^/t����y�B�N����߫Hݧ���n4n(��bH��ϫ�Q��O���>����ظS�Ygʅ��g��WiN����t,�
Sf�e����M,7R�]�ۀ��܈��v��)<"T�AC��W����IM;_���G�[T^1
a5@ ���R��<���'k(�6��\<t�C�nv�7z� �,�"�����S�Q�"�I�:� N�����#��=e�H��(ۅ<X�i ^<���4k:E��nuh���)����t�tR��L(���C��cEO�����LW<7���h��ۼ��"�s.�o+Faf�C����/�fT'�r��ׯ��d�TOD�./��4�ZL2������erfv��5u�L���pK�zCǰ��#B[��s�گ6�β��y����-M���Q���. ��p`��2&$�^�.��$>+gݥ����1*DLU|sK<QL����H�!i��(�O�ݣn�/�r+���������NM� ˖�έ7�р8�3qg�^���=��*�&  72�+�0������h�&�
�_�)�$_�&n�	]V9T�F���Q��?xп��(����Q�0͜��Nj(���:�>���S˼�7m����T�5����XR3�W���6�X�d�q
��XmI�6D�"F*�S�Nî�t�O.��uoS�Cǉѷ�F`��S��
WF��+��l.tE�[�����W�ې<~���P篕n�e��	�gO�b�����o5�x���#6�˻��LoH��\fUle��MiR1TrPV!��4�.��1Iw���@�!�R?��&�#�@d�V�$�1i�U�<�ad�N�q�s1KiP�����#�Բߋ�n��_Se������f���I4C�!i�Mw`��	�rc<���.Lҵ��ɖ������HϞ������p�X�\���q!D�k��o�Ir���'&����~�z2Z���7l}6f ��IBrn�qo:���A��BL��%�R�^mH�����2�2���^/���,�(ۘ�ѻ��m��㴀���j�R(�}�qKh�"��dtgn��0�d�/G֢��P	S�l�_�O��Yg�9�Ptv 5yC#d�ɭ{O
?�[�x'�0�����ӡQF`�0�O�YV_�:��{�t���]�J�{�n�O^/�	wͶ�ev�w�I��S�o�Ң�N�<�i]/��@!.��̀	L���
m�z�'y]S\H�k��N�E��v�mq�x�1F��t� ��C�`J�a���l���$:K���?$x�oӶ2�d��u�R ��7���T׺/S������p��'��{ڥ�*e�f+eh������rp�~��Bg�a��r�Z򛳗ʟ�k]Jr_���`� (9<.>�%�bވ�����[`Q;�1����GO��=r`+����U��(�hI ϑ��iVW*�3��߭��������[�nl^�+�юv1&q�;%���W_�#ӕ����I%���V� �a7�w�u������ң=-�E�J,����ޑJ�ȋњ�z��|S�t_���;��dX.6R�A�-�Z�V���M\�h'#���"GdeA��ܩ� ��
G�v_r��x��K��ؕ�P�8�t�@�Rᯇ�|����u�d5�ZRO}{�����~��>0A��Cv�~��s�ό�㻼��Q�^����{����a�>����p`°�kR��[���r��{>ǘ�C��b���"b�<�QG�?�"��Nh7rh���$c���^���g�\��lC�B>���_=^�P0X|l
������2�hȖ���Z���Vqŕ�2��mQ��B�� �,O�cv3=�'[�ӶW�e�0}��3i��4�|��m��0:gM`ǋ<�D7|��}�}31�[7��o�2��,���4ZȬ�`�7�>�����0\�2Ioc�Kb
�D�Q�L���:�c�����e�yO�G������0~�u (��M���G�W�8����ɵ���m�B����]#��X>njꡠ&�_��t�TP^ߨ�v9�z.�n_�a��{�%>����=���T�VD԰���x���6eP覀_[�lJȿ:�CR�H�B����M/��������6z�m��P>���W0[�p���E����
=@�y�����CV���Y/Pt�gi�vicz�K�8n��HC=��{+��~�K���(h�Le�4o�-|AJ^3�AHf��P��]R�ȟ0�Z��5�����M��W
�\�ѿ�܎;�7�{�����ZD�������==�]�%��ߝ� w�o�������d~Cfa��
2�����؜���AH�綽>?�n�9Ǜ��\�T?�@������K�ې3��[H}���iR�e�WuMQ�6ބ��X�/;��$)�B��J��mwU���e
�0�.����3�_ƶ�IW�� h�����h�M*�n����U�������*c�j*��.kB���ϥ!61�MP��� �;���pC:��F�lH������Q��vͺg<Ȍ��*	���ÙK_�r:R3�W���w�UT��03/�.����-c�#N�,:��[�_���]��W��/Tx�g�v�" ��f�l�>��`�@�_�����w�؛ں\���_�4h���F��-����W�A����|�@����)
��A�R�j.�X����&R  <Ȉ��L2]/���h��y���S������o��mM�Z�_LH,������-s��LQ5g,����	��%~jc/�P6>�Q��?���m�` "����R�Q�>	��j�����v��qʶ	+�-%�ZANyX�G���\��<i'��->"	��o�גuu� zު�=��~���\k�b�����>�RŔ�2`�;+����4�^=}����8u���Y�Gua��QZz������@~�$��}��Gr�"(����@�MCp�}&�ȉ����X5���mX�kʟ��]��з��Xs��/�S��t�)Z��ڈ=�h�jj�0E��u��%���r ��M}w��-0����n�!ecԥ�j��h���9�4-kIA��/Eg�J�ܣ���J�Ilru�-ѕ�ԩ�8IN�c�����F��:�v{`�QW�0n���A�ƓUJ�}��1.+y�iF����*�]�rү>E_��	����xꬬ�H�Z�W%6�i��õ���Y��'	f�I�9�;P>�b&f�q7'ۑC.�>Qfz�m�Y.<���x�|.�}��*y���.��i5��[i6ǹ��_�24�^��	g�t�?1bV|�e	?oE��'�98̕��4G-�F��\*/
v�[뾪Jc�-�T�e�ُ@T��6>>Nv��EAљp�E3�5�����>n�7H
�JF�@NVߴ-�?��앭��bt�HL�Z���h��Ƕ!�d�����6e���F���|E�����i���)UbGK�d����#�Pj���ͬ�>�:�����ߜA`&jP&�V����D�����\��̣�4	��j�o�����j��P�F�C�*�zH��x�d����#YE�f�L�J~֭�\�:�.�}�7l�{=�Rg�T%wڐ�y���qbͪ#΅X���ʣJ�������!����o�|�ҤD{�@/|,�5��l��bN0�ڠ��x �ŏ��xJ*���I(�������g�Hw3	����Qa�y ��H����~�'�m߇��z;�2��[0	6k�S��	�9&�D>�t�!�~-3w<�>S��afy"�5�o�Kf�ҽ-/�.�T%�wځT6w�B���b��%SF���h~�����ZnoDr��!N�`Qb�-a���_��Hg�u�Dm"��%?����s�,D٭h�&8�Lo:i��{���=O�.p��i�b3��J�D�Ҏ�V�X�ȧ�G�v�}h���:�����cEVYfP�-J~X��E�^H����Y���V�?>/eB���5�3v�?�p���vo��ٗ\�#@�8�f� d����P��!�����L�	3��Cv��RFo�*��F��1��\�mӽ���4d9�
��T�j��a_o���WJ������T�����ƺ�WO��g�<��@~�\���[��W���VQ(�D3P�F.;�F��kq8`�C�s���%�)���'���������m��Y7Eu�&�Z?y�ٯ�v��	�����:R���=���Z��eP��}&����LZ?{�5�Y�+IS���P�&��K��%q4���1�H8~8����"}	�ɗ-Y�p�io[��q��C�q�d�P[��Z�ؼִ� �W#P���[貝��ϓ�݇����Q���@f��$U���0�V��LA������8��fH�7��E����QюR,9��Τڣ��ds�<��-���>�7C;�
�Ѕ��8����;�"d���Z�s���Bm�D�'�	r;L�IOWZUi��(�ʡR�ͺ����H�EC���L��?G.���Hr?Ӳ��t5M��q�U���¤�����N&c?�܎F����r�����G��m<"��
��X�/�r���^�ٿ3���#�����ʝvw�p��O���G}l�{��ťt�WtC츦&�Q���PfnNs�C�� ۓg,���5�� ީ+�ڟ���]�f�����±�&N���U��OJ�wǀ��,c��Zd��� M菕*�|� o�8w�����߮� ��
%��IiZ���ޓ�垳�5��n	���(-(D�af��ǈ�w/�v������`��K(\�й�$SëZ9��3Lū�RGI�Gr4�AH����Q��6	��1Xc_B[��z-$-�/<����*��_���j)(�Hd����4��R���u���	���8閝7fC�c��|�O,fu��@����8��	һW�^�%����mWU8����a���=�֪�z8�03�o�>�G' ��M�g�՝��N����LG}�dp� �B|` �d�ߡ�,�xp{N��fu��5�!J�OO��Po�o�S@��zP&c2W�Z)���a��7��ɸ�r�,Eve��W��bҞl��W���v�!&�S�,��E�F�v!�7�ݨms4;��u�pF��|���dW5�50|臿��%yL�=��?�\��
S��{����t";LX	�*ړ�z3v9e�<L���d��aM9㚌L'���:DE��?M�wZ��OV��k��*��<�v�yWB����q�S�뷿k<N�B={BF͂��l�7	�`�kIm�;�:6��Ȭ6��Ƀvq~�iQw� g�o@B������eJ{�%�G��Y�%1�A�M��,����t4р����K��~�ü���y=�6��j���*�K�M��B�q����Q��v��sh�Ӥ�YP����F[���)K-,������0��:�PU5  T�W&��v9"�;�f����aV��F���0Si���5� 7C�C䣔(�e��A-�������]f�KUUQ}#�<%Э`�jNh�,��pL�/|��$a���վIefsW#�]���%T6Ŏ�O��p������ɇ��;��������oz���q��j�i���=�S�`:��/)1>�G�0�{�e0����[�Ѯ���(c��������\΄P΂uoP Ξ��b�Jc ��d��]!� �:� �mv���es͵
 ��Ae��o��b�s8�k��{!��L0���%���qi+�"�(L��$����5*d����%���ִ�v�Z�>~Ǡ���Z%�-!�z�����h<o��g��t���Zщ� �^2�`����T�wђ�]G����×������ib����_=A-��s�4�ǲ��9�'�4�2e�	H�� �m�� �Z�^V���Z&��q.�\p�쟕B�UW)k�xm��}~3�Ҹ��l\��=2�W(�����!��ʒ�����H6v�g�pZ�tF����)	�m��D�'��Jp�;�̑��&�˞iP ����ޯq:�sb���z�0�C�C��/����l�}��F�٬���U~:��e��u-��	\A"6��B�ӬQ�N=%(WN�~\f���\;��A��]pՑ.R�7���n�3�.�f�����sk��+^�RT��ޮ[`0���z���o��R�_B�2H����w�od��dAs���p�:�r��Inc2q�9��
�ch��F��bK��x?�tAP����" �GL0#"99�jI���Tl2�`�j5�3�G�_9�aM�����zC�@s�]��Q�Y�����H��e-g��e�\���ѥ&LQ|���	uѕ�-AEײaV�["'�R���J-��4���T`kd�$�XsH����Y��fm��Jmo� �?���c��c���������׌ҋ5���x���g ��0-_���M׀!h�����-��Wi�rm_̍}�ĳb�2bؒ��!�&[������驂��&�r�.�N>�a{[2�\�yi��(�a6,�
���1���w�`�P��d��zpX� �3����9�|e8;'bv|F�HM�{l}(�MA�?pI&��g��B!1��{�S{=���1�_�C�Q{0m\�*ĂH�4lE]a�GA]�_�oop]��&�ԋ�X.��c�3v���CK���k��ϋ�Q!M���j�C����RJB"��j�� �u)C��cLaל�ݲ�5n�;eϑQ�$)H΁;qB[Ԕ{~�X�v&��q> U:v��?�
<�q<lnc�`;3I�̱�˴�w~�V�Z4�x�Q���h�@�ٮ~Q����Z�G?R������ʂ��Ø�R��i ���U��yW�	R����F�9�gʃ�����x���Q|gόʛ��62�3��Е1s��o~���A��Yʓ�Dv�e�{�^2a��$l��7C�2Y�]f�8�:���)���h[yꖥ�6����`!��X=�1�F)p�Ҿ��+��+����!�J���59Dx�m"�T�DY��>��<.�XO�{�Hj��jG��='q셃��[hq�3����7�kx�=��Yb��؛O��t��閐�m&�U%nE���M5�ar�n'����~̾&���M������U]�=#u$؄���$I�dw�n���jHYBW&b�W�)�M�o�����b��/���h�P�~�8!8a!���1�_Y��B&��.�F�q���et>Rwݔzz�?:(�˦"��0�L���o�D��4j�6�Z^r�7z'���#��h�:1l���\iGUq��2�f�����6���\�f]�a����m_OR�Nwa��1�U�/ƫ���Cb�q5g�1�ƅr�Ĭ�F�O Ův�Sa��
g����f�g?���DZ�k�z�����.�x�e����(E!U�&lJ`e�uM�0�Mҟ�/���A�=�U�����V�}�Xi�A,^H����9�41!O{��d�
C�k�:�sp���Y~��v7tb�j��f�g���!<N|�l�a4����I�� �Z��]c�RSTp��� ��W�fڪ,0��m��訠5��B�4�s����vG"�Zu�E���e"�$�b�rM�ɗ҈��s�čR�]!�/�~C�J���+�a=Oϖ�?�<e�� b#��=?cϜ=6ⲭ�ؘgC���Q�*׸.�ₔ��5�/Kpǆ�P;�ِOWXP�%(����C�ll�F�A+�E�~��C�9}��_mi��/]ua{(�$6R@L}ق:j`j�}YH�}��Z��}��(
ik����W����}C:���%v|��c|(���-#�������E��_�lɠ��z���܅�gy��	��p���e����X7\�%IC.� O��y��d�/�v��nj�>��	�u��� ����-��w@؝�(��}�2�3���Zj:/+���Hi�R�N;�Kx��Ɓu�e�o����W��<�A��h�z�7r�:/������3`�E]�T��*w�N�gat�\|��c���J������G��������N ODRQn0k��������&�U���m���>��q
BY�g�"(>�\<ía�җ���"���̂���ԋ����^���U�B^QX��3�qAJŦk���+��[���^�:�[FdŢ�o�:;����R��3�8m�DGܱ"����c�"+�����OF�h�Q9��4W���$ɇ���Z�����W/7�8�g�CǏ[T��*�JGx���y��2���F�c���V���