��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k��ib#�Y��&UA��?��?�%|A��͟ĩ�x�Yrl��睇�Z�Ǎ���M+�|҃��4��6��1��O�%����D=�ߝ$�i�b,$��hk��|�FI�w:�
m��:um��q���K4�a��^T�6<�q��2�ŀ$�����:Qy����o���Z��0W��_�V㮽28ߍPU(������$���6&�6v�g>��Nw|��º1�-�Ϡ���jS!�S�.��� �������6��UY��Q�����5+Z��j�!?���8�݃��p_���o���ZO~oK�(���ʚW^#q�p�=0@����y�ȴs�N)XX�r��[��vld����Q�1�X�=gQ>I�i�#��"5�j8�;&4�ŋA^���*~6x�d���@��U��n46R�Z��x��Q��{ty������yܩ�N���T�G�3G���4��_�\ٵ d*~/K���E
R�5�v(� E���^�y���C���`�@y��ci���������g�E�mՁ�{�H�a{����͇KF�C���W�O��e��8� iJξ�_xĆ׶>N� �ۏ�� �	c�'nT<�s�D$���!w��#�%�k-Nߵ�="�U�-�q�ʡǷMε��Aѧ��QV҂B�6D%7�M�|]	�M*2�<~<�n)}������&u�x�daՉ��i���ɐX��L�E�J]��������܄�����r�ze~�^��l���g�����-yKH��d@�
��m%	>�����+������������:��L��$>{ƺ�1���m��h����M���}(0r��L�)����#*���v�/�hM��8���'X�����_�nlPN��z����J�i�x�?���ҿ��I���b|b1UP*?����S��w�Ww����߷�u���b*i{k-[ �!��&nzl��Iwͩ+ZbZ����r�Hl����'V��OvmdWi��Co�,|�U׺3���N�(�6C��%biGTC:6�;-�	�1[&�]�����"pOHyr[Mj5�:����'�A_Ė���h���G"J6����HNF����)r�d3A�g�(F�������tpA)}�=>��0;~��I;���FҔ�$� �(�: j�� �Idx��Qb�ϩ?�^���|n@Ov���[����rK����K�*�v�胗\rڽ-�?�]�ѯٓ��\�ZP�A������M�g`�4t���ca�/*\�)�j��!#� ��������E�aU�O+�~�^i���s<�\�<�_!n'���YV�h���~����٧�_��ѥs}t��%j���C5bS'8^x&��<S�A���$H7nG�<���э\���s9�)]!I��'9���W�MP|��ɼ��&*׀$�!�ۄ����
�q��ٍ|�im}
$�n���|2O�bU��M��Z������S����Nf��v��ٮ �:�Fc� G�[^��ɦ� �kć'<2���=!�.��w_6�Hm훯�{��9� ��b>�*���
��r]Lƚ^g.R��ilb�)��D>�������D��x�W�>Z�ɮ�!d[A)z�y+�	H.#x�©ͼ7��)9o�)�<V���Շ#��Q�����ryn�-��u�;�~��s��J����91p�m�V�W8ަS����W���à�&�1��Rh�Sϊ���sb�gO���5ZkehaIW���<84��@�@!Eh\�Ў���Z��+�X`iO��zh	3��l�f59�ϗ���:�z;Z	
�:���A�a��G�Bk���xz���9��AAx�T�&t:Z��xd��si�ʗ���4��(���J:��>�@��S\�ѓ���?�UBe��1s�Κ5�ᐺ�.a�
�~m����	��L�)��u�}qX��	B)�6�<��ȅs�m76�;}���^w��^�´��Ia�N�����v3I�D��$��0��A�>��%�L��Сo��l�g����F%�i���Tn�;rGWJ�3s��V����ZmX�{���z"���K�r�n�a��Ƃ��}�vkװ%�c��[��.lb�NS�%ҁ��G$c��?�Da�%�%��>E�H�nV4>��3U�#�%hzd͞�v*�%^ء���U��b:� p���}�C"U7ǁ��i�¹�A�C��,��]ų<�J#@"�j�����z�2g,�w�~���O��n!��t�18�7y��Q�Ċ����\8��Q4ü�f���f
��=���٦��!��[�=�ܨ	ط�����Nނk^ne��yA�	,����G���X?��RMx-^C��CY�/H
�#i+,��1"p�Dn9r^�U��CtF<'� ��+�
M�R�n�H��d>R�P�ا���c8�=t��S��������s�s+7"-s��W4�O�fp]��&!c�^*���Ԕo<k���PݒPR��zx��N��}|z�ͥ'uRM.��j=M��'DI��\rИ尿���&[�n(���@"@ދ����㆕c/��~`��RL���A��=��x�f��qZ�V�Ǐ�?�AK �'}�`a�ύ�s�Wf���5�^���#F����5�K/SG��b,��6İڱs��gO�EqZG��<'��[&�.�D�ؙL|ѝK�R�p�tD�����A(���G܇��muMc_�	�Ӟ���G��B�J�ߌ�����pEY�����=�
���ce�$���2���2|T.O��r�[����mX�[�~�Z�e-��;�"M取ųT�+)�Ҽܻ��?,���R=�a�^?k9i��3$@w�U|�s��9��a��	r��]^["�J��b�!M�IvCgٻ� �v�W![�g }؇g�;�	k@F�D%LEo	�Y� �uI.nv^�x�E}�}�GKGq�ah7J���l��x(�}-�֨;�|�	�Q��Y-�$J�����D��<��vt <�X����X9��'�ڏ��2�R_��k��f5Q�V����o`9���s1G%n4W���V��A���hxrC��5O	;.!�^5��R$K�襯�%�t���c�4���xÝLK�"�����J9����(p�훯��o������{�x#p�)8��!?�����a��^*o�WU_�Qn}e~��"b�e�l����{�xH�.<_���e|��/\?톆���,㷑�y�YuY?�x��fADnվ�⬁�q��6�X�y;,���3��Da���L�!�BZ֑�4�φj����}oL��F�f*6�?�O��=��G�p��GX3�\/L�K<Ou_�]���{E��f7���