-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AScJM4mRMMmelawHT4OwOdjttUDOrCJVAACsflpO3J3nX+e8z4Y0yXST0YTTs9NRac3Gf6vODgk+
R+BSX66gXn3Ly7zsFw6dOGu5T00B+0U3nJ+TxkYtDhPCh1fclvDFp8FRN2aK8CKKVeEg3Nr9sMAH
k4w8GsKTXnFf8iosHiFVWZ9Pi+V9NTLM+vvXPAqnhvNH1nWjWLiz9XBFID9KYcUnK0oaf5qhY8rz
TcWGL06EOPk3rTc098lNtUQTdQyA+GgMvuxk7+AoY46JxHgdNcP6Xsz1QmfS9gQOagXvtLkksyip
wcQbOYVeFWyufa1p4Jh2BEc+iQvsH+zSY8JjRg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
hlDSgZp7+zq3TxHshCIB3o9OKMKQ0B2r+pWcSM8kTVuhA4BVbzzAgvhgVcMZHXkPO/dxEH6CDMQ9
J/istUvNpZflwPa76G0hSVd21jlYltGmFPib6XMq3I8Q8pTTu8vrPr8cVjZZSpXTlj8MUWgS9dE6
VufduTK1uKpPb7rNwm0ikkN/Py7eCKnI+qfVizUbgyHoukffZ7WnLEupxJFZydKIvHg6S6h6qfoJ
tAhvSoqOJt7rWfh+DqtLTVSAXf9TzGuLzHk05V3Diwp78tSH3A3/AE8GAJxZ79YUVgQlJK3jrdDM
UIVEntKc+pVO2fHcaVb5GRaHYbnCIxDIZoAg45tt16ZAF67qcnfhj+u86a9EqXa6HNhDC72k7fBW
z5RWa/DAZL4rQ7N4rauclc/zkuO0ffVXGHZdycCND8w/w37z/JerO74RrO6oN/EBVNU95oSFPLeX
tN0ZNZZqZGl4ETs2Ljp9DD7GxDdJSYpm2Kx0IsVhGuC/fdGiIVIHBOAEuBe9iwTM5VSGO0kSkeuL
Zg95kxqMsdRdrUTpiYBhuzr8CsyjyuBI/tIlEVFmp7AxdcsiDYFrt5oKD+Skrh6Kc2D2G7aEqMd5
XNBOPX/wrMDEq9PY36OrV2GCXcpdkBKofSLS7gpL2EKdl3FVsDGT77MRUwZ6gUv2HM1RzQMjRdiz
uQhwb0SJvOoi55R6dfpnhHCqHEYihZ8VyiB/IuLmMOuGqcD2Xg0XE4wnZ77Y2r4JOP1Nl0G12Haj
A3W7Rva9NMRQAG5s111GXcJTo9OnRQ/Z4X52gpT3RMa69f6YKZp+wFzf+2l8ufAvZPJucQ1dH93J
6oVrzgGZ73sBW8+DFIsg0pVw1Es/F6+4Zqtfj+oS+eqRWZUzSn+kWWGUL2mhwsljt0JAIxrWhB09
0FQVUYH0o9XlfhRgkNaAxPaqKlUBecBtfZSjX3gbkI9JxHDe4dOIIXrd088sqXJurtTxiCORM0gt
lKdiBWkKqTnpofQkhJl2zexwWGzCyXllhoac5th/KS24aE/9dHws5QGr5uDg9co3OYcy+bvLZuId
f1dHkYLP2N62/1mW/EcGWi3vntFeoIbrnvIMt3j8p82oF0QYQ0zTk/GHyaLPBk1619kvrbPHGfX3
3iw8kFm6OzxYM3OvWJLNTbvWHJX32QTyo6eWTB/smCg+B4PgbzoNu53qxgxFFRt9CxuQLBh1HH4F
33qkVTCHr1bQr4HDj4P802l+Ksb75dozs6zLNeLoGXo/tmIm0NsJCtKS23lPVHEu8DeLk4g6c4Hk
7mb+wiCInduKAkiJfF/19imXIIouJ1TYjxfq6TmxuDf396LG1bMNDvkV9vEMkURA0jU3DgBc3CVB
p4Hp/Ls2iclRP6Yqhfy0nqoP0U+WPa5UITJgM3Rvx3+8MX5Eu3SEp60aTBl4y5+KbmBBldvSoq7A
y6s44Y8XUILcXqEWi7htJH0uHlWQskMiYLllLR6RXu671R7c5gB4QukgvXnljC7G9ObQ3MtDZHba
Q65EZnNdCztZ9RYvQnbNyt5IVjJahwRGFXiqRIURb7ROGeFhmHEcf2+hzqyjV1HkFUuXe6OPKp0u
l9+wYAFpjH+0ockoICHOK8F6BuTPK6ILXMc5e59pY/JW9fFlqmoxGKwKyh4n1VggFmI8VG/F5cfn
7aPR8DF+FvfnlVVzSwaewwnJDweZqIg9LaBNZY2MGQYZwRgcZTMexsLkFn34cZwPfwZ5JjrAuXls
eWqUCYk9PNTTxP3xeiXf0rcPil2Nllrshh9JN3yNuV25gwJe18AtnsSBmwfyYgIfL3kYc7bhXlMN
QUNoJCUB5Tp3XAevsSCkmVJtirhkDpkogDjjOT/96G8eDPhb1gekO5faVcRGFpJjxVRWsngYiR8d
FUFCl2EnTxX1C35QQZQI4d9zfK3IU9y41PsxaGhXWgVwUmkRMMIo8s3G1/j2QHSqkrdn86/yF70K
cI3Lno0JDJc3Bbi5zftSYVvvW3z9PBtWah5q+bdhty1FXaEJwm09fojOVo2d1atpf7PmF9PnNUdc
XvWxWG1tvRmUiiiYHokQ4FM4F8LlGX+UEXemEMQarzPJgWz5Y/qiY32en7VmkOp/NGEeYhg1bD8m
ppbiKVElBwPJHLzd30ZIWvXT89nVqzcqov56klJOnEWp5wXD4gygBNmbsBVwyI9JjZ+xiRcZNXac
I8bAKMMOpDrD9ZsMd4wKUFinqzoREzoxagXmD7AYMzXBkL2AzWSvMmpm3hd38zrqhIJbh7M0JVzJ
+Kb0fDzHjkuCpPYDzSD8JrHM7gXE1BLkxUyUaKzifMlqvOMsnSnjMPmde4AFwdTExDVOhXWmr8a8
fLRdO/vksfkAUhe3K2POq2ZJqLUY1NpWcS3ybJ2RHHSXRzVoT8/RNajlSKpES4QwleI+jV+1YPqG
elv7JQnPLZbKs2YxWsW8rsWFyBtiqyt4/vLOnJ3ivLralUKq61SCnW+vxooU/45Btfy/1RTL08S9
5gGTlpbhA1AEyEc8vBdUSYAWI9OzVMZ4EYveOVPzv67JTqE4XkHlFaL97o5BtGXLfpJCLnv2x0Ii
9yWeUiMjg0exeRuCm9NVDqid+LrIMp5UP3s593MAT0JvpWPnsqRvqMzD67Av5R+OVJKXEsg6V1lX
vJoaZ3zcHX0CiUfAC14Mbd4q5kl38rI2G3pNp1Fh6oPIhx0Q3JPDP6EvvlH1/qw6W+WXe451NiKe
v/wFOEWCtyKbyNfspBkhr7Iz8gHG/kV4hmUgNFwrAvqKNr6p5q/LO6FCI5xwwyCj9dWQuU9TWhiR
AuM12Mm4hp0JqLtPRD4ip/lwvg2vTp+Pz9Ym7C9StwspSs1ggXg7klom4zMINIO8YJtGExDQMO9B
CaFTnT38EcYsh2UXCQcdp5LzL+stwkNQAhdKHedcLxrhy7dAHRmRotTEVmMgTFxpf2K2MH+db5m0
cMszIuXm3uo7EXXN0GCax3DuKMq5taolEOXVPgyElLCX4ZyNJlrmj749Ih6gpc/zCMw/fF6sMSOC
ntkPFlrLD5xZ+rzdHjdWpkC8xaSgjftYdB31ulRnNACAsJcboLbrKI/WrUQHtorrM1r13DYZSXdd
CTCBQsCzdil9t4ebl5Z33WBewqnH6E/B62FK1O+cj1oV4wmsxRWZoDmIG2Y5g1rhyy7UB+Ne1Wwj
oOgu8nwk/V9ww2HRkH7XBqxwv3r8f9Pk9SOY4qMjXz3fMymiDShcpRvyMbJxCi8RokoMQaYBYldN
5pXg0xNbsdsRIeHda1KRPUvc9R2q1/FhXybuzZdzVPFYV/P0DooKGwL0TJZBj3XWKq8n0dYWt4HK
dBMKnmOMFYcaLpwtjHqe2L97w/DIfOt8sLeWyW3zuR920M4wJnOjEHUxMKe8UG4tVpgZ2dOl5sqk
Cot/RDHfmkO/Z7rznT3kTcCQWXKANaL2ei6Fvk8NOhm4swuGReP9Yv+QJ0+BjEm+LED+ZMZhQwOq
H3aTCHn6q4KBFb2kc8pMEMSxPK4O2/xndzaoS/CzPFecQXscsuOgBKCsG4th4v3zcgFnJIO9eLld
0UHJ4X/Rq60oNYN1zNbDI/8e+blFlT4a2tRjUE10JT3Mvi9GH+2NjWf2cz3FKz8ZfKvJgWV5aOkA
NHEMo/iRGINZbYJtku7U690zPNvup4zpg76nJoSpVKQW0peYWIkVo6qeiU1VjQFSxYU2Eb/lx5QD
ytmBt4TQD1ps8MVUjEQywdeCq6O1dJM6ljqlMhcHqg6H79geYNr32IGFj/+24MDzKWpKzOQ24xr/
NkAiUMDUjNfJhRXHY/3MI1uLEC9OYM2srU6GSLxhq1yYTjErYrHuloGkvClfYTMT247Ltm02pJ7k
YSXXb+Bxs5d81jan2UFLJfQnvTalblmHGMWBcKOgQLck8/5Z1oyfl8Ovp/stzg5TtqZLM2gfOFws
XV58GbL7mFfW+/Fmii6tJJqICpuiJ3rB00SvhRweEcB6xiGxoPkEgKMKoTgZFi5wiXia01CoyOh/
Lwpi52c6oifBmTVFWKLZFPSmRXEUEEmyxiNGNLtsoxww5gEQuH5Yy0wDXn24jQ7NrKH8PWSrQt2g
uC/1lvlrkt2T6WXhC8iF+5KdQWRl9brM5SinjpDUgRQ/ytnjNIg1eESGq319XIN8NdRekZBnbRTp
/qiETccC1suuPoltdvxPlpnXBek0IgbchlBytbdc2++4Xb8Eek0EovHTEkC2XLz/DcpsHNWJaAmd
y6LgHhsq5NtnaD8iZcZV8dDYAEY5ctzpjLvybxQyGGP3ZWnRAvByF1g4cBtq0BsCfNNc8hAgtmOV
ylBcw98w4PlXMDOKLmM21zGPTggjUtY/E8Bqv8YokPF5rkAsd4aVA2R8MTE4cKcItLgX/JjErbyi
Ku/ZZMqK1DtuXUSapYd4//r73Zg200PR8R9EBuws4spguXJ/4NOAnOPUuRuKs95gUsxFrd6lbXEQ
QKqJ4JC+vx6XojndJ2QKc4oAoCPW4a4LbvRDq1CeLSmfNjxXwfEj3CE7VOLdE95L73tj0Y7K7K2G
63DE43gkmrOXTTed9yJ8kMRh1lOGYBl42GdHHlK8Vl7QdGOZbe+z9MwsRMaFC7DoveMinaTPRKco
SxdFRkc8i6TG2LODN9mIDvEkHAeoLS800zLk1cJf4nkU9kceAt9Kf0XWg6tRDD6elog2jXIz621W
2Jp1OshSnAgJPeLFqQy6/gWvOU5vlF2K1+ls/MBcdONjATDNybgfhn7sm9t3cWtnJkDlVQbBqXiZ
0uiHAU8ZrOsnaPq2wU38NUWkloF/Rp0BJDD/ExFhQyZXEW6pPVETisU7vqa7KvFgQt3BZw1s843P
q241UefQJDqUUA3o9eRlU1I57vUw36q2NfKJ1KJ5CtRIqnCTgyU40teMzy8zjExpP42tYKuLnm6X
ud84nU96Z9JshHSpo6HgT4Ti7PPdS9zaIzx8UuKU7p12ESKB79OcSwRA9cZeb5JPh6Z3VinYyy9+
v+t6mQCuVysIUg9KM6ZJ+q7lQSYWIfgVQroHJfKjQpsQ8NMG1B2j0FDmSlOVa7H4s9reT9SHjoEM
hv8OxWhmACl/IFHxvcOjubezBNLrloyscM7drtTlEaQwCiPDWlB/SV5xRhpT9m4MpNw1/2hUTydc
OrSQKo0HDESQyWdB9Ut1H329PuXVk8zW6b36vJWLdi4PDUWawRzbuKX2Ecf/2dvTKkfInZT7Uoa9
V+EXRXhWg8kEtB7Sr54ReKt9F7PFtPZAp9QO2Iz5sdVNOhG7LwlOJ5ocy/67SHzCDuUNzEvoZQwA
Peg+geapH0Rwpfl7T2AEMhAUy7B8akMAhCAA+Ne4f3kIY/tIP2KhaXF8/bM7k9fRX31RuphVNn16
TgOvmzSOuvHjp9hQlcX88mIaK3yQ/aKkvwD85ivCXifI+Vva4Ipyc/8JT9AKEBsVqdy1n6aPgI1O
osJyDryBw3uP9ZGcEwSy6g8yHuW7dfgsfoOKUNmmPCBJ43CJt5iWdAIp7m0y4sES0lEykW8i5XMF
bJoBQzqHc6UMylMa4CBP8KhIZbjsQ5LYN04+6b4VwoRHS2TzEkR4NCxBf82R8pXcKMU4XTnwkVby
NE70rw1J/1CtSGuYeyoMPpnuo29DwheDt34NaTbZWlaEi8nYKIg3AWHbPDfsB+weFC0tKRkRmnpN
5C4SoAuRI4Wv9n9UBv2FzNk0BaYkJI8eAK8uD/CPja+VBEPy937vr7kEahVbLBIZNrFuKTqnH7d9
3uY6FQi+xzIRzoIRtyIBQs1WuhaPNWu/YO+CIpKeRs2biMQmMUVUWeebrf7C6/g5ledQhNyUXwCz
0Tm1SfsEB6AF0rxE76kF3DjWWNEcbKdd+QxuujyURLfXlLjuwb9KpMplzXDD3LAFttXUyYErR1pW
zvL5Lgmm/yf4jiuodtdcjabmIW6mxELnURgqxYP901f8MWwqb+u6WJSedFc9ZxvvkeirjfH3N+rH
Og6URdXR9bPOaLGryJ4ycW0cjto9DytuvqrptD1+6jEYxXrfqJhxcQoCOLt7jfxMAoaP0HryQSMe
tYCG4xnermBDgaY8G4h+g0ppeiTN08gXQR3PMZMcU9SAgPnsXHFLrU4OsZR8ZuFDr3ZWILnmiytg
aflcl5DzMQ/S8/RjWn5XCk5XarCjmYhL0EPMnQoS+gYUkSIa+iDzy87qnfmpN4phnVgAE1nMj3oq
DwzpmnOcXgcBjT5M2gYcQ/eYsUINK555PM8WR6O91e+t2PJKREQtYhyioJTiwDUtx+iRVqCpzds2
Dxy+uDoQTl3H3TwIBdm0BLc5Qg7GZDIcM+Ahkv6gCV05Fqr2I9iEusKCZaEQQYKndYqbK7Dy+DS+
k2OEagyG0jK2rwUdgyNgiOcvAk24BxloyDsEH739hSj/NCL6lMljmT9UXTQanEcoQ2xuYIKmTtUg
lhL4TEWat9DLu9wAmr25Dtewv1okVjL+F1jSgn0MgcqFc0d+6X/z1f85pYQS1n/2b2cl6Sl+AZfQ
GLEVPmovbW1znvcentA9MPzoDiAOMFNMjeB9oSmWhgvQ9+wGcllvWnfnGI3U/7oruGRXe8XxYyOQ
Pie3ln7kDJDj8uBklWCYSGGAqVNz/PxUJPgTOIFi3vAW1YII5KOxEfxciG4n1A+5kqOFSTDKvZ+2
kQO5jZPYr5VUbRkVpmK+ZnZ1vN2DsZIQN0D1Klg0o2wWCK7GV8eYruCBD67qPTfnny7rq4NQQcdS
YYyceut3UCuygEqxbO8fvET7FsYlcQPvos/wnn/9R/mjtdbgJ4E75GjlWAhFie1zUc+3pkLEf73q
5wXSWQcM5zYHRJ94/POEgToJVt6r7TQfAjSE13CKYUYqSCHCsJQp/NgAQTsSo05z5vaoKUG62FIH
c5Q4s96i11W9C7K0hR+MTcfl5HINmCEV8VALfOed5JhdWmy0lF94mDE+sc/n5cRS2KPXylPqn+aI
wPdpOATRzuv+5Q36qP5ssR+zWuubcaqOfDFCs0c2jeSXGz5lEAbuK7yZDBDKpQdmcGFc8KV6XUAI
TqGHXBuraz+N/vpB7ctMRrMw9l4QTnXlRJ0vi29DJtp9Sn1eBoe4xrJSVQYOrLYazYHj45L0iZw2
pxYoSbwvepf//BoGLYS9VnMwh56Lemk67lQJ2RpSdKq4Sv5xlodCTr+sqGCfqSAB4TMLriwA0HL1
+dIDVgFfiB4KjopJUxELDZ5zlGJGVSBotipGi5jmtLypPToYT4ZL0SZBiiIENwDldIiTT8wiTksA
S215347/eNGATRKqcdzNisi4T49XYbF7xGMZ3RyQZQVeUPsXM+qslrF05F3BKExUHC9JJHOiiQye
9UfkgukqMJMpsbP5OKNtcs9DkPJleGofJuZIUnHb6xjxKW/y2aJ6Akpz62vzKIlmfjcuz5773KL4
eNiMu8kCAMiuprabmlL4QI+bjewfiKlDHr7B+uEF6A6JAMPv0VCYJ0mUTKsxEmZfuvE7g4Jj4zxF
lt8f0ZEp5SEo+PL2FrgseeTPsgjygZ/TKxC26MFrjayvzXtDOKwZBYjoskf1brt9nxNAgRhzAQ+E
KZV8E0nIeWeiyrribNzwe4v+Tnn5LjV7hxUM/SY/dYyIXqQrBHrIDKQyht6UkVDev2NWOm6eHXDh
5K0YNfXe/3scpdVDf+mB87nZI9KqQ5NtKhnGmMkQxH0j38hvFut2y9QTO6eYYWwjilWXASFJwJv6
eL+fYZckv+eBC+SsEh8tuZvjoLbaSfTm7olT8a8opfab1h8DNu5ZGJbd8rjEorXkN/b7wlXa5J7y
ZkPrcA4yCA/y63zZbzvYKVd/ObxUobM3g7F4b+OHkmDlXYwlITHXnrPpap9htQcmRghZTp1kOit+
8O36TUx5+FrmT78D8VEv5s8oLjd774xo1rcxgjzEFETtSA25dx3qpWk7brbyBZYRzp+0pcmosESW
3ufleIkxvqN4za1917IFq5qJksxdDpOp56QESrJPg/oqPr9Q4oHUn0te86x/d3FCp3E1Hf1ek+Kn
GavuDq20dFyO5rYL2FRccxMgpNGy0oV3OaYeOt8e63qRlnfwCa5sarwzOXSQkiwwjzZYulco7Vdc
Vm6poPNtjZqeDPruVywlNWB6Q3IDWKXto8Yy0Ol4f9flE99Br+GN3bZSw9FmR6QmLChepsbnDEhV
ATJhTHwR0ExRm6SRi11mWRfomSxXv0+J0Bxk4oYOA9sIVLTJIM2E0EhDUTKdM7JZXD051CD51Fsj
xmp+cicihkWulV/OE3BeJDLLpVQ5nBhYREc7ESJuN+Y51Bin1oDJgkQaS+wgVWlT2UXPGUF4iWPg
HFT4M9ovv/XS8Lpc4c/d5cy9nkJ5/UuUA1LNl0TJW2UDF56xAaSgoIRXz8JkWiK9wnz1B/FwpXXJ
l55ROH8mcRzAbtOSgCwxyJ8SbKMqR9Nnd7JjWF6pxtQFDde1IRy8BeqkSQBxu4zxbccn9iDEe8+9
0Qtvx8RClYypU48573HzbYJY9drb/VhXc510OwnMX/4hwnCgYzAGXJT2BUxro8fQO/hJYOJDxL8Y
mymcGmzG0wl7xLKih3sv36YOKxym/B0toE1bMZEudJ+vpbtF1W27xqnPg8I3VsyBXY/sW0Oy51R9
MvbEUazOVYhD4egKLKFoCAzyBh8zO8rpBsjCld+XQQNvPsxXaar/VccnY4w2ZFqDpGJj7mJerRqx
4qKdf4S0rW6gIf5DjaF3IJvINz1PNQn8n2YzKjx0B2fBdPC06hPB9Z0hMjVfBe6liaCKgc+btuT7
HXKYD/bAiuXcj6qZ76Hha2KcZDvSJR5uFG+pmQpAcEeMhUXIqlj37nrlJu2/t91wGSm0Ig54QSKn
Tiv3ifFw3fXCx9qbLFJPPNczduaoT8uvuzMCtc51bTtUhsYQndaXDf3VUyls0OtNDcVYNQbd2fBf
FgKXNend+YnZtEDzX4FrKVOJZINJKfvtXG1xUFen8Li133sD6AsCU18rQ3pWHsMjUFk6zj63ELVs
l3EhVgqTCq32BOqQK4olKZbcjRNfpbYTbwXORZXSjkFBh9aRYVvRXTnh9DbQ9/vEfX3adrpktVCp
+uvAtMYoPC48rmucWRQt6n5Q/EH3a/qJbj1JonvoukWo5Wfqi54qxDhfVeSBbnDWdIEXaz0DZOOU
fPey7t5ngEDDkFFvANh+05fGFa6sMitfabpUXp4/iwBtN4nx1SLznxl4TjkhP9t0ITGTQ6N7Gej8
FkRoV5yMD5OOOLjWGZ/KSyg0Nk9yA4pv2dU8OtZMAJtQWxE5hYOgOaswIlj/CmAOhH/qCZuAZNYJ
DhuE8oBfDHZXQ54khXIZ5HH5gfqFGAchxYVUETN7dEGC/iqxWplAHag/nTUQnxUJT72PQMWfQZWj
OvH7y9I/tgu0E81658rVLvT8AYki3lo0qcfizNHSkIbZrwszRNBUDD5N1OGx1nCTU2psBPY2TpN+
3MR6zsLnJ8zPPSxUDphdYk0n6weyVdxS8fuRZ4XnccE7vQPuDGVNoA2nqidaOKv6ekfiDKWWdC1c
CLzdQHwQmo5Z5TsmQbBebWCf16cBaBCtEz7op1NSyGTSbsN+qokOps5BwO9cJY8YsF9JMrCbrTbE
Yoe/t3exwtvqljrKXhCnTlr27plQ6rMaAIB9jVgc6on1rljTNp76z/UYC29ZAWkdwN4wbPoUqpII
3ZKNytO8xaG7NiBk8trmFbrjlVIxtqgy0H0FJ9X1wufPTH3UhAM+azq5+J/MpCXiBXKhBOlYjkUY
dv+Q/zrDP4WHindU89h4Fon5MZZJN3olgVbxY5Hd7eq4oS+xgZXwXqtvIEttGyRf8flCf7F4GFs1
zFkd4a9C7ACJ/cDZYURTjXZiNdEvlZGkyF0E3IrNFZf+8aSYHlI18ixX5HnKLuO7mEjeSqa8bfma
yxpyAXjXHVm7Nwx2lvDkNsQcqPOVFFNJUncsh/EsY6mmNWe3LxxBKJi0P0YqvBo83rqD6dkTdw4a
S+B5r2vT2llqRA1TywM4kaG8yFecelypZQ9HmrBGStnQvNH67fDH+toMl7s6RpkHrqtHRSvLpy4K
WPNCo0myBZjhmBs64ljgxrL3jUTux3/GjKKI7dHaau9USBtIoVFYk3rcvLmXAH77xf9DpAtfp5bn
XZym3W0te77n1RYqsgSo3bEC4TduA90ZFhvSjOOyoJf66WkSjXoxBVtN2pJ+TATcpK9zSeN7n67W
rdNV0Se8tN5oY+Gf5bRO4aYxst66Qdsl8ZhC3h605L9ZZ6NJFxcUCFRRz4gE/XIcJYcwEGnZHtRX
/H1eqZMWZwCGEZwCxcDDX+PrUeMPZF18qyHemGWhpi0IJLiEbLqE4runVQi5AltZnZ3+5De2fH4v
HYj2aDX4QYQkRGrGDQCYcyWzb5KTZwDG169m5NktbaEmI9TAbNfCN6ZCD+ZyqNyZVR3ltsb786EU
1LNwMBOvMyIJtMPu1WqhQPoMDyk7u6LhAvKPnh3VKkbDZczjx3dtfB9BReR4UQtanXVxA7wlWRs5
0t1VQzluuwupxMoHukv+G3GOJoEu81eHtLUCqh8QfvEhrOta2TyWPk1oogDcBOPaDzSje+uYAwJC
gFIq1DB0f2rHhfjboUZW3N3ZbPVmlRS5zRrdr4amPOeiTrG2pncmeP+Tes2KY+4l00ojF7C9YvRv
1gyC9+oq5hBKz1f3jl2la2zNCCYcAPrM8SsdZyiMQkpZFnKRfAlSkbz3fhj0nMDhqN++5MSG0Dtd
tREHVgz82/bzw7q6TIl5W9azVfITj9Y2jCKrob4+tKhrfAU2BXnZbH7fvJwpeXHWrUxckqYHTOoy
+/Tv6OyOGJL5fVwAsxNObyreNS2v609cCs3j6AfmPfBRegMAIfFKNzvfd/VLykAZq1mrfRulncms
ZPEf78hjC0YsOFsGnGcvrYbpQ8cs5VanzaXWz1J9bE+xKsKmRmWPCmd5DxmjUaCtEpq4BGmIeqLi
jr/qIDEM+OL48GM2n4ZFri6ijOO+iCUfb4UGPV4ZjbrEEf7+4DNAqNwk5VOplnlW61eeb/ooT4yV
xdGQOprvTarNAVKLNjv5Lfdm3CPYAQe14uKSmXD+9gKgHRIkA5lCIjVODXTYcPwQFBx5kxCoZTIj
eStnTVJcNgiK5KBcUNnQeKIlOOkdrPsRpE9VsZlNcA8zQikyr9EuBfBvcDum+fC3HyakUUIW+D90
hjLMRnXewhMGvpGJauBnK2uXYPoiTKuqjdCe02hcC8giJ9z7ap45qCawk/KZ++KE+qW90Hx0Rdmq
BJJSF9vERWLQIT1GtOHq/8X2VTSHYsPtzea8oBbof5OuHXNYFzjregV9BIMe2qffgLMmGso6QNCd
lAkJdB9bmFUEjspCu6R1JkmOQVvMavPWLZhnvSdrVYIMubNhAeXCeOmfeNl83A09N5CBDqbYEMi0
cgUjfKN1zuXd/UWUrMiS838wNszWAbQB4fiD/CUAllIR+5rbS1xb9d1kqiTVBRG57l2M2rwQc9Ze
0PyNEpjSjFqjCxHRF+7ozr9DE1k3Rzow34qdnbwYTv890vdmFpOmJgOkK8tPs6fR4sC7OTaAFFj4
LMiweKI7UcS0izxdF/tU9ERQimsjYObp+Zbssm5w0E/1kgfy00nLH+eQYamizmMDwbYzigXu1S92
l7EYomYax2ua8KqjmalBfKJhSRBvUdESOlA3mBhCWpPfRWHMDVEcKwpbw1SsdGm79KsQxZciuZRg
J//ZDHy51C4hc2rap5SZnBVYZooE6Ui5xUqRK/R9Z4sTK0KusoK1rfhylnT2tJLJ4bg9tw6FB68f
Jp33o1tqV8dDALaoq9iWidAK/C/f/+FALQzzHYhKqw7qgi6PydACSelH/d175YHjO9kWgoYEZ5oI
67zWTI+C2UsJj/AWWjWCSK1uzRAfpG/J7saWulBOmCoRqCIxEC/wIqswyRHSBnUTpLJJhYEmrFBv
Czcmks4CQiwI54H52D3LnKDOxyARn7gILDmCduhsE/5FEagXLHedaehKc33qogTuvHbjJEiMCKb0
Y+RyyNKszPz34p86vojnEazGOI6nmPNpyzKWCuVQIIYrm/N5Zh+UYdUJ8iB39fcwEahsBjXmocb/
g5l5uKQigxZLzUhFiXDrhl9pdWXFR5bxwtY+o4Xr/7SnZQoAJD3Ih3Tq3kBVbLwI+Asod86r42fe
YnppT6elroiqg3RROAK0jKODIysjOUCb5FaJTJAsUHbF9yTaqCb83Tm6p0fLs+eXp5niHHNej6Xx
r04DBSgzZnycI4gLfXv6im0ZRq33+gRCcyLzkZ5NOikMYy5IwafS7WG7iJyyLdLO0LLPiP9uvqd7
a8EcrcbwSt/SKyRyNwAgnnBdHyBY5QE6rXX2OcfM0pYZEA+b+5ZyeUivhbu0kEk8mTJ2CyeaBsHp
Q45OTc2s6gAqnAjTlJUqRyhCf7f+OUs2zY07Cefk8m1bvz+EmSqi6h6rDBLuwUaBRwvv7FBraWcA
iN2YSF2wX7npAjeNy0JJA1EKYuEX8FYbtmozTDtpnHMo2LpkjtLiwpsw7u5JSMUVDO+soP0rh90E
lvcbIw1MdgLNKLJTPv0deQG5638ZkZnYZNRuJWqGBUQl/TZUd/clEqXw7ti6OuC+u23gAPh9YwLA
W1W4LkmMLkPO0yBJpuss4oPBdGgR29+oqQHzcfMoF2dO6e9DNSnTCY+nsvsQiOPX3H7D5QP04eEN
2GM+K09zmUfFuojwNyxCBhfUzmYhm2Y0pL1XGQ1VJ4ETOgpObxjOG5mxbuUsbyJRQIu3OamJ79vl
n2QTKEFO7aE4YAI0EH6X4yN7TN4oZ3JIznLTaekDeN1FG/j4cEowkeu89mbmBkjaKnFO+7ScT5SI
q9YqvSSr4t9LL0p3T+TnReaGxNWBN3WF/t5JyqsNcGGJ60dqMmPe3BrKFBoKhRtJVfhe7HfQlY9P
CpWsn0HKgwmGPsWcLg0ibCEHnxqhYjsY2vyHGMAA7T76W1uYgBtYGPCu1ANqU2NBAuCaS177SCVG
8w3L1tbzD5/6ReddINi5KQn50kSpzCfLV6BUgyCBV7LJwQ6V06neDJjXvoq4CoMwgESvHJNIRvJ8
ajsQ+mzJ38ABTj082XHWElc5DO16eCdDq/GSPU+awesTD3CqjiPh80ium6B0okqPTnj2X1ZjGCxr
5LrB1PS73hF41wbG+2ZS4rnF2unfaBXlzi3UbezTT2h1nNzkLQP4wNZ1FNOeBiB+A+rsuZaGbaUc
xDfXbS/5LVAPvQNiG/N7PETTT/SRY7raLJ2Syn2N4CXA62aSGfUgPpxekuzPLJwOiUL3+do7gIwd
+3y10Vb83P8LGVHG2lM2Fc7VsQBAZH22eByiQV6aKfDTmPFgb0FlFj35dkAB9mX0hDEArcSV/KA2
ZIRzKEZcSoD2d/L5kyw7Te12hI3hXNCQG9FgTTmdyUMMqPJx7gdkRw5OoewRrFi+sE5A/Ub1klyP
dMFbPgWaf9shvWpyaL/izIYNCTetNonccCnc9mZzUt55CU9Xi1KoFzo8DAzD5ryLsagcRz95DoCE
oVpelBpzVEoX28p37NtOY0QVpra4Tvm4n8RtEJfpk9YaDYHYeSw0aQqaaNaxte4kvmFnAMFNY+0C
Gt5WHkn3t2XZTsag4zlBTtSrTuy/zkdcHVat+eP+uoja0a0EBocxwOGkJxWyTkb17nWhFUZc7IA0
nYNidNxwQBJ0ZyhuQMhr4ZsPK7KvVuh7s20tdpQ/BnzXAjY3G/QQ5L8wK61mkom7IHcx20PTQPn7
V/T9ylScWv0ELXWp1Z2buwQd6IbjWqgNq5KQtC1rjk20LefI5fetydVuqs+CgdkIFPK1r/T7axgI
lSsFgboJ56b6Jji459x9khDFkIMa4erlhoN+abX1Z7XsW6R/kn9BoWlasMAI/4UW12RI6I+ifzaW
7074BSOel/BjwoAe+woZU2yO0NBNrQcWhUzFnZil6E7DWvuDryg2XsLbuGnlGMxCUS2kwXJ9QU8B
rJ5sOZF8DKXByu1AIFrQ/8Zzr77nHDihlKFNWEfsNzx9KeLa41OEpN9gsswzc6PuBWm7CbZoBVhp
m3uf6yVQWTMoszcPCz4DGWA9AqkVB53FTXtkprL2+Q4SCsMWRWYReifLyk4XQJCRQjixY54aMN2P
wLWDUrAWl8X2u/2TPhlX+lY1EvYCwBMrdkbKrw53nKQ441UOYfLkMRAcTiFqH0e2VET69ztwy3yM
kTTkcV+YXRssalurGLb8q17+ZtuoVYK0n2j2p0Kj1ia6qYOv/+5pmz+SZzBfQFmWctQCZxppPfXk
WiAKFe/DzUbtWa4LVL9LObTfDC+IOqlp5EfLO6FbJLhpoTndQ36FltLQDKzoRJkD0L3HOfV8uAai
+hT/K/omTvVM61E/DF0pME4jUpTFG8ZOSuHfrL1zk7ILZcKxrTvFzC9NSrOI/Q4nyRtTxwidRjS/
zBCJuYFC6NEywA8R+NqbA2puH7R4tLW6peAbqT8bnE6DbSSoN1ZvK7FpU/M8tRFEAlJodZsOPLTr
jZoIHdMjk9cOoPR3XFH8oMfT4DqpXF0Ez6pS8yK+Y86uNkCLM30G1axnXatoklV//XwLuDGELjwu
JMSxKDGzugYNNy7hK4GJfBo56m/j9Kk4Am3I5TdjaBthPhPr217jvZa9kpQH8Ib/d+CVE0Ol1I/J
UE4B88AJJsbMPzSz+MEtQu36F1ZMc6mjlbWCkNiDVKpkqd1Fz3VeF9YIqPnNdeFy+S8bwksvBKcm
L9vyNIHX3ysgZsT6pXnXcOnS7YBZB0nzQVNJP+GNLd4XK7+4NFTgGTUn/zIVN2jyKRePlyeWR+cW
dAjVdw3I5+2hv1YUgGSDZDMbKD6AZAItJb1LWxGd0geb7gqF4hSzxdeY6GRpuYs2DA6PtEvAZ7Qi
I0slSehvdjqVx1VKr2ziBXn5yJ0Jh8s1uoYEAc/h7tVHo1p2JWPNE+mA/JACbctRfBZTw6CzqzJU
wwYM6Y/jbW3ScS75U6PziMLZkF+20Wz9CDgUe6coeClEFHt2UPrvGOw1hAvqc41avMnbvNfqxwws
ry+gWmU4bq7d6L/i99wv1gzqvF3S/IJFcrZvaWZmQTwo0HD/s2+V7fakssYT5xL7i2x1Tqu5T2vW
+o7zEt6Pp8Dqm0SMMpW6pKl3ll6VwdtjJmffSwWuK+6hwzExuhJ0L4fkzG6a8mWIZ27/iCWVtYFS
JBUwAkUNE2WAWIolvoFckrE0JDkGu+9uh/XpSw6iDtKaLmU1sJ6RbTzn803Y+x0kMp/fLBfFlh9G
4ZVxsr7SeuT5wgCOjk9pQh5J5CIzMWFWxK8fz3IpG2HnTrXCmJwTsZ3eMR2Fhfh9usQUA9mrbSLH
yH6y+2CGf3p7L7aIT624GjABwhvgUnRmrgzcJkotwrJVllJuFkvNSF4pASnkZMIMH2C004Jc/M56
yE0QCtscJap0W46d4Y3NNdTPRwLxfxlT/6dolBm39gAz3sUAEVQXm7kCI0bgSI2NInFn+B2ibzaJ
3y1ZDhXAgIjHlFXPqHcnvrr4z1Pydavlq91QbnYzTraV13r54ONyrCgqvfgKQqF/GWqGl81hXB1v
F8cuU04WxFI1CkOLMhk9YTlhmm1cA1EjUtWJujaX+1RVQW4PrRhgwlKvwFve59URzY0MoKLWfgE3
pb5afD3+yZtxRpUfZw/ohuL12vUg3222D6wsPwyClybUVP/kffMGsevtaq/JHKGxgdSyFNXqc/k9
Wh1oq8L1OfCwMJYHJoT643frLfRrhfOvWQm9ckmdMa4BLawnJ3Tu0fLe0yN5yEkoVwJ9FJxuv2Oh
fFfrA7hlRQ0tZPm6HQyxc4RkvPRNjLdH1o6mFXvLxCPU1QQ8gy8zawnRUUL/CDZHA+ldE3Of9V+Q
juYCQlzEosafVhewco0FyJdoQWTt9XX7K66of6Nsagfh7bEaWG44/Bix1WUmZHyregBTpj+R5p62
7V09BXnRwhG/f+afa15alFafdQEFOlqizwQujqxAydxO3OdNXo6mg+AYVyIyz/5/wS+3w2kinXts
MIquLK/L686POa02VYidqEwZXoNtw5b/LwadkM6urpDhYIUc5MneqoeH8XHvWiztoI9lgEANRePb
bSBAj3ey0JvtMEXJaAQMNO6kn4frvQdV4rceRWQBfyb1Re4RBjeMKdp1IHnPWjh+uawjk0cNLLxc
6M3RLrwRxDJYxXXHxudTT/1wOzeU2ObQw8QebpYEmSAG8RoGM1nism42iuIWaYaMgFwmKOWFEMuU
QGMvq0+wTtabNhLIHpnUX9VaGlgmdOSxhPSnx29FoyUw0GoMrWjl+aluf3ediyjP87neeM94zH1p
6U7oLh3eDVJbOYSHMMeRhYb0gHtiLgT2K5WYIpOfWNZzxQC2kWO/c/Ocp6bukNRWZagYzibZr104
PGc74a6Ecw5Jvbf7OZF1mH0+LxRpCjfELe78ZYKdOH12MBviJKc7KuIfAJISR5Prie2Ex3qeZhLV
89tEIZbcZwUs+MX+ACzDSspKItUTPPQcscHlAWVSisRMw+WHVW/XZOzXA7CcVt0daWm0n50HJnBt
/6yOhTJMlv7npnuzeOo/FyASS5fqQb+l0xLV9r40RurrduBOh8aLSkIi3VJZhWDfxiU12yskcF49
MQ6N4r3PdaqNxJbgarpDRwNm3DWHGm1UDDv/Xa4iI3sAr6+eA/oHtqJY1sqAbcxza7dJWx1AKwRb
ogiIDZKa4zhi4W2Q4d5a7J/uionIq+ps2C7uPh/yX2epETiFlUiE1sQ1MYemDUKofUbUP3+OP9B6
RuYEr4WmdKTGwfw1t4ARCHRGkV/uMJ+Q2yAYEHo2pZ9X+Y0t5TuuQUe+8kr4SM6S/Q1uHFMj1ehj
PNSjp2QEkGUAdClbnJkXsX/Mhxc2ohqf2JHt2Jzgi6eS41z0Cs3HsbafG//hp53Fv7ZHglWXnxC1
wDeXFjC/CZiOa1Gs94ZR5Lu43pvK2d/ENmpmH/gXh5UF1lBv1zkfogjTA7EyKdCsQGDpKzSFU57L
U1sag/akQNiOb4FLx/dNWvumuRXA7e844XgSDHBw1MSuDj9AfzckTrZdWk6Xutrz/79tjbqzWcEi
2bw4Cb2BzUl+wbt7CnXEae52BxUkwOj0Yi7UjGM+sWAgN+0QVGvQ/2QFl8q9ex1fA4DnfjHLJuZ8
KypOXV/odOryudkK4LXnLbx9rJmurhQ35WVQRmKoi04vCFDGXM/Jf5eGCbhY9FZFHW4HSAV95ylb
XyyQ1y0wQjZQ77oVHhyMabrNR4eY0E60HG1y+yEExH+0U/j6KSylwdhIe6k1O0k7W3ZFTFcyDNjT
DxkMYOkLcuLK7fO+rWePCRNuLUgW27SccaVg+LuHbFdJhq2fVig4irHWepjqu9dJWHwzBKBzLCy9
NWwv+Cs+D8RgMuqPCY2dtBrpexDKeEyQV+3whkhIbasHVYbjVENXf/0ujKAmY96noivarv84evbO
qMIViAt1Qgkcui/AsZR+eF4bxGHZcXxWnEU8hJ5VPfTivk39ekjBoPb+Ki23qtvVvXkkAPCs36Dh
iNA8eQkMkAXkYcA9tDymOtYdm577rtmcliqY/RZqSfqwFVGbv+HjhTuuRHZVtasd0eD1wAop/Mec
UEmKiDe6E/w+5JAWPvntMxEC2KFD+8ZrK1YejI5YkAlyhrVdP/swfrtlYrqBteB6aJZhr519aI8d
zu6DwpTWRbo2O/8Wt6WCNklIrWi6zYamJvjEgQdmLyK2JMsPmCmC3xq90Nx1TlocigXaX3ucDaI7
1XqHfexufScZUU2vN3HrG0Ij1jxAFD8x+uNneH/ql7kS+KqDXEGdrgpgETcMC9Wf1oJfB4aFKubx
LnMdaRx/MeSJdq5l6JN9Z9rcYOvyP6vyy8t4jiyF+Lb9tBa+LTgD74ON9LIEl0iX1XJkPhVtjEi8
ltPeFMcaVSnwdGErT3cR/e+E+eQmFz3g1lCVh9K+ZB1fXH6RwBo45+Os00iWvM/XMchfg5p7xsdb
vVcL30QkHwRSwXhq8xLxj6yN9gelAOyViQljCro1jKiQFgloSEcXjAnyKLC96FJV5juZ9to4qwnq
olYHrYFYAMxduF61T0B0UFrWw2XomIdiZE6b4fBmqQpgQNagPiT3vpeLjxqXWfS/unxpcp4YP/ZR
/gYrwjBLN8/UlnaaORXiAGLdubeWoigr0/U1jLRBvMYWEw/aKltvLfaNs5cqRhNRGfjfF9kqEyTP
jMdtSenP6mAgesx7lIjOUPT8iiR/ZRI+X35AiDsjqxRzuQyKsrR7UrTUmTWaPwzIIeJKUy6uK6ei
Wi+gX1PptseQD5AtmAfXPBhJwpGaeRCb7+Gn9bpVpcEyd4xnWOmTYHPIcE+Kc5K95ZADnBIao0WA
xwBxdXq5VRHOroA+ZHvIAk8BNUzfgtDdA6X5DItz74PpPTyiwTVsyuQORUvrPN4/22qV5JmYB+a/
AnJzRahDcJfdNJf33dg32KLj0TiRSIxA8ZF7d5utuFzuEx+qpSI4QyRGMfg5IbONrfJQ6ttJG2OC
3aVM9aziBKsRaFFW24WhOSpt0dH2zfbbI3915Q2a0GC+1fkqaU87/rXZ5HGq40GkqMxr6TftgBk6
3qyoD6NHjQgvErFBf6joZmyM/+eRq3XJPKpgnX/En7G7/U48JBClKArbMxf4EDbnC4hsNoIwcGgr
FtO6NNAc71qUEhNBupJTcJS4/Vqk4xGsjdimMJnY2MY+J9bEtwV6SPgNDN7JiAVoI5MjKJTuFRKw
r5PzUohOBO+lG1qetBb2kUUQnEjgJctDekFGo2O70nDoMrSaUW8HbBSlO4UHlt98lpcaX3l6o1o0
3nQPu5BmFe+U3QXn64V7g96e67Riu/8xBvivOfrNJOt8TOiDHjVppFZbnWbnzDMmTN0FoAMN+6Vb
Az5S1BDdFyNfOrPhvXmNI93enwSLyzrM1WDsyyZQdAEIHiRPwFO41hiBjSHSliHzzE/Fj9xoCedR
Ry4cUAGlxezltN/l5HNfXE9B7akNaWlX4UfHy8bmPt/mwpD9XkU+M+DloKwYkoAQx0WADkluw6oP
0+bREFGA8vyxF5njQDYrLGysxD3AyomgyCi+ObjcMooGsBXJRdKwlatbxsmS5Qec8xBSQQBJugge
qetgXs2vYMncR/L11v6StZOHlGxcFRlmHznlC2Dz3YRUNvI7EGOuX4ehmY9NKhGNnH3dHQIDLeOd
Ox605mbN56v7fLOuJt8ee40ZtH6mMKx42GTRpp1/brhJDci2enDlp5MZJtlI6SSXGDDq5pQ3f8Lf
Hz3OW309gKwmxunzKKKbHoq4qpMgNSab4VzSexvg77OiHpuRnDxVnEWX16Z4FRfBMiUHhITkJzph
us4kR8k+LGoXkr+r1seJ8bnIWBb/lSLCsT+NrJLQecrvp7KORyOip5G0MERYvBPV0OjqaXlWow5J
TfBJ7O936GjYOfJ5dNgKuaXRvrCgY3uGpRF8kGm713tLwZHoaxmNFDf3gw6Do9fkGav5oBKLr4se
tWORaXl8IfQ6W9QwuAgnLVAHhItieq1mMpEfdcFDE3NFJJJTJyRkV14iRAdoVJhMCUIzkGjvmmQ2
rFAySCR12txxowFk0kovkL1rYjVm3IsCgge5yB5sGNmA+9Sl2TQ/oCUi7nNVjl1UL1IUQy49vd+q
NhL4Crq2rDX2TRB7YepT+3OEK6Fl8AZFbfZ0z7LrZyR9gXcE+/xltqtF7qXGQ6rqSmKSTVjvZId5
31L2IgUK1gU+GqVz8mMUuK+3t2xDuBgtzUIiaZeAOCLttdJHYUSXABBWfFAnbbPhYL3xjpOTX2sV
dZY7EluScwGbrIpuIVoIwm3bJ4WV38WE+cZ71g12fpRmZVruGULco5LcKxmthlfWOCsL/naiIP1f
4TRJ0Obj8pSUAh3yn0Urp/x9Vl2LPJJgiWdYKTUlt8wlISKLngBnmJY9gQM9snbRYbtoyccgdqKb
EJpRj8T2650x/KjlzNf6G83k2ZxIzpOBcf+ZKj203++JiIwUboqOYPz+TEVGgqTBVPl3B1no3PMV
Mh5VUgmIGJ/+nRLkoC6E9+BVRdB6Iw9zRaX4sWx8/fuLA4uFHMbSZlVXtYyy+CSyXJoHc5VLBHW7
UbK3i5SjmHeGwh2gDslcKzRssGNK+FNQi6/ZOUD2oBwIPqYNoB5zN00SEtptK8PbaB2f44noBYqa
0xcFcfWUiJwizihcPmheAOWpCkCJKFn5dHeHCt63wXcdJmgb0QfksA2dsEfX+NwMW9iFCdKj6pna
/YRlXyhvtAhK8ZAXrGJItGaITCtNCvedf8Qu3XkYUdyO7dPKsEv4w3EUDBxPNhISlCrnUJe3/Agx
ro1kMF01npqt3zEwOg6ETYLzgkXshNwv/yx9ZZ8bXZt0qKr+tFD6qeX+4dvJ1/ium54O5+8pLDPW
aZPDDJj+zTtV40pb3krB8jTWCB/DgnqyHps+L+24UPajDZhsqNsO12x0oKSZWhStxaZKvjdEv58R
Y4+o3FeZceNpxpa0thg9+Iqam1cj0WcAtQSwZVMRBwTIGiYGEmxa29jwuycP+6t3eie5Aj1wVE1W
5ph7+dEz7yaUDpJcgIYSzWcH/MlnutyBwwZERacxi/ZvNqxi/RzzNEmRYyyh5ROPy7KvyjbMKz+s
AGCJdUPrRXQsgnBQq0JFUFO+v6jzs6pma/bFa4SOeGJBDxC9F6QTNGzAFk4aP8x3+X136SYqJF61
fu0i3bCxW6mMzU1FynjQ8nNGhMteDI2znSAtaSI1Z4ahTA8cZIlZd5t9zFIcKdnxhgICCJFqIB4s
yM+EDk9vLg/tG7YPGV7kdTquqVJNvl9Qf1mgyV46lnNu1Et1efJknWpPpDqIZJ13haEvAdF/ABsV
O62uJmH6OgleiJVwDP14sh7Lwf1kskrymNlpHNW83fPq5OUU01EQwz12U2WaurtOka9mwQ+OfT+q
JKd5xtHyz9QiY/DgwHCjDaKlK65WIcZ3iw1yGAnJ8t+zU4uFM3Qo1mpqFs2w1nFnoAeflReSYp3B
EtyJ28Eq1zF66OzEn79oNVyeEobQ+LxW+HW7UsZZn4d0jLpMe7Qhi+uHQoEHInxg2z8DQtX7vi0x
/UOxjhnr75iCWhH4GB0RuyO/Kt4EK/uLw1Qu5XCV8nOxOOZNyyRLNc7TczJSxE2Ky3AQZJE63CvR
NvT/6XQIDSjtF0CdKsV35lEY+C3XuFSlppGKvCqIY5ZwpSlMYIuYERCcz3ucAp+g66BBi7gZiQqE
mINvAkCqTaGtEOsedrpc8UHF3BBLCh8QCGrfDsJOMBd8g2tVE7Cq/g7cyXi1p6UImTSY7236s0cx
VsDNM+K653VHq3W6RZ37VdDFtL/JkBnSPYpKOt3r73VDqvDOW+3IVDC/KBSdLa8vapzt6g8E5Uf+
AKlnkh8WPYADNQry4jMAiCUcBCd82LJG0gtujQuoZdLtwSu9wix0SsjZL3Q/oy7q7EAMD0c1Gdfq
vuwZ78GyK//TwvXjG8rd1Xeg/E5++SDF8TO2CWPGUPDErGD8DNie8PFlxbOIZjn6PbPSJEnrfNhx
4ZPYipFyUCIyi/Oby7x81bo6/ldh7s2ar64cV+OEJzFReltUsFq3fvRMRZw1Wk7cGb+XOckcHuky
2zznzfBp/SVGqz2pcn1Y5Xz3qx6kKijuK9tHVIlc/H7VYNPP/AMdoakLAspkA507ChsOPb3Ekvx0
S14iIllM0M1m4OBteFX1k45wba0uP6pXLpSUfwUItSyKfAylBvXeK6bFuToTmDl7m5gWaf5bi2nr
Yo9oGQ+BZJzJgFZuGd4Jq4XNDXMSBogKN92RQ++hy6DJJ7DTcLQR2Ho17HkGSvVuNbvF8iCavRSb
4/lUboa+ldTvettKuhQRvf9/wADDCWLNX/jRjWfKjSFNgvnz1DGdiaCybPyIvuh0Ib1fFeGFShHM
gVA55A6x46EjPWkEsPxrpEoMw1MFXHv48apceyqV9IZRKRqCf0s5KQxlF6Vb2RUwWCz0Uh8idGyG
sgeJCz/qAbzuqRIL43m9CIcogMz2rNQXK0D2s+EaNHqRVrKOO/S4+KH5GDVz/fnAvtFwYbvEXkTY
gc4BJA+vyA01WTA41zgDvthHeCV38vPTiIWc7PL5aiilpzjrJlbm8vu5gSZtfh76ljuskTaoiaGr
Y2Cb3IqRm5lWSJUKJAsSGLxSVBOTEuqLpx66JTsF49nJTK61FHVjCkTvBXzVu+tPGf0NcIcfFozb
ATtQIzYIWf95h9edDU4iwiOfLj85EZAiZdD1rnzC6IpKUFmtu+2WfPeg+t3Qnf2ZK9f1MGO9HEpF
aJeK6TCotJS2PB82iHT25vKcSovi5rfLxcOkHubJuIwmm6ZPyresXHDYvKQLoKD2K1F7rhsFcMPg
HxZrVf68D7O+tcsHJPu4LU6p8TAHbGzdpGKDD/XKY1ZJT2BZwYGs5HY7YNAszCiKZ7SYW2hTiHg7
cDPiiM4uSItTgqvq2VnC7zUGaGThM+UIsGU2u6C+stZQ4kRs/tXpYL8e+87FIoobbKywrrzkkc8V
4XXhoOPJp3CdgOgWLTW2aJyOCqxZH+3bBI0nOoozWDC0Man428IXcjpzSDsOuHuwQ1+1qIRu0f/C
wu1dfrNyOHwZ+36YZ3tjOLyurFwU7h3nti9tSCOXbPuurRtL2beP+/wEi/fVi/OkWJOF4OI6YYNo
oZ/IyCx5Qa80YahaXvGuO68MB6iraQFKeA3HjV9k/HgKq+duAQ3WybD3BvZXrQDNMKY/BWyasfBC
Aq8UW3dSyTFE180A+TvVBl2sJUJRJ8LbDmEOMnk7CGKMChM/wyZeRsrBtBtSDtsauSGUfejZxBYs
hDQ0pCzSZvHowAfbe//g/3TL4Ad1uJG7RmeZdTmpCaY2EyIPwmQkY+h7avdrGMrvKfqR1fEpVNjl
Y4J+MCbXULfIEWuIen0ANNZM3lAdcGhg3KJjAxxgzvey0KeA86Y4TvqaujSLO0yCbBJHEHC4S/V1
4zPZ4QX/x/nIdtSW5lMjAlgx0wknY1f+Jv1KW49dYWUcg5y3Khi6eAjgYmfcbSQIsdAky645YY7L
JfCt+I29+4m2Ot5h2P8nQzRQmLWw7zCmXRF9Lgka6SqP7JOFd6YQJJxGJCnl6/RawnvqFjvq1Eph
bf8bA+ueHKYz3NGDbSVMT8E7+7CcaJorP/MnU5dTU669+o8+hGkNtMWWvXAP8zep67MFALasW5b1
Q/IWaGreFrliYkV0OS0714TCV7O1alN6JCCM5peygM32LoaZJ+dpLQYEYxEzzrRumImbyZsGVl4g
JSSmPbO97J2fzDAU3IQGb6XsUtaOWW66cWS5t6zaWLL8TRmVYMqLwT08OBUdFfZtEQlt53+1ja6L
cngm5F0V/la4NAovmfUuJ/DR8a5QDc3/rRjFE33XgSUKXNfo1Gx+fjDF+MGr3rfQzjD/779B/6t0
1SfmLN+ekqCBsgVwoYMdB1RFKpe6zYmF14B3wt4J+cm0oAOAWUCCRHJRug549lOiUarE1Pzrj93k
pH1gyrZJQDoVfdU2Fv4RmTWWSQjJBCvcVhzh941pjR3yhq80TnI96hsXjBm1Z8M/P8HidO1pf5Fo
yqihxGZGiwtrZQ9yoxr5WOF8BHPkFu3fuLR/C1Abj29dauTaQCAEwbV9+PLGjBEEK+sDrdBRrcGt
WwzZowMUBsM2UmImnvl/+3TvQl3RG+FuP098zNdzx/wtsX0aCJBXC/1tZWvCH2I4+0YiUZT5MaoF
J7w+38g/IfelhqKt0A1MOpf9Q2Lsfpebj6THnhRMRASGgvedqLG7Z2quV9afZPXI5K5vUPJRN8Kz
njegSUvi6pldRWgwNC7PxNJTv5dIrdb01dKUepatf7Z0lp6qqVKayP9JnQTyzj4GkUfA8SV1LgW/
/TImb1qI2JzVDNBV8/8k/y/3WzWPThhCirG3SawN01DmtwE4Y/45nOYZB30Mz4bUuvun1+mty3gQ
1GBCZTLFwoeezdWQcPpd0ZBd2VLoLYfSXaVYd+A1WE1eaMwoZNGpuWIoEFA6Cgmj6FwXDlT5yxss
6XzFE2//i4wz5hqvgPONhrE4wpLPDRnivlEmGsMe173kLR1H2Wd5V7FFdzY/Tav6w9kHlkluUv8B
e4YT5psw6w1sQzYVUFUfybvCAXEcIc/9BqS+eGq48FOxfJpFDAu2vwoQRcBBK8NuHUE/FbSOZeem
WxVld4flR4B72P/CmqdJ18AxIIKpE3p2jHRyOmCDjuidZSZmdvrjDSdK1Fkzryp1KJa2LXDbC5oF
RoXj6jAvc3SK0VCCWSCzPz3ZDb0hGFNhZqAIDfo8VqsSyqIkqwmercRGK4zh1+m6cVQqqK9eXjWo
H+2ucCSaVtee6IKC6pc9wk5ThXkX2uu6t5EnYI0M7OKuA83dK6CNp4Loexu8lF5E5teknUmpE+PO
cv5WLah0aFG3Hln2soQnS9O3ufsQGMhWFxeFRBJnhNPgfjkIBkoZilEv21RPVS32wD24BTeiZqBD
8SGru+yOx10hFBmpjjpLPiIyjh4NsxG5bfBAechzVqf5r1O8VaMMO7qJf5JhBT3VjeNunUaWz8RV
tlbapdm3MghdM1ouhsbJ2a4rPI9LmARyVdtog9zcOlp80gyLZYvJSQubhc0urMzv+scajb8v8543
pNeJwl/QRUDYMXPhwRao08oJ4EBOR5dSEs3Zxf2HGUJ8PuIvhT9imLTsxJOT5INg5qwTHIPhzGOs
OxeElmlXzUWyp304uWRkZs6+z8mhWZwxbOoconble9m7tsvqpcEoiVKfCBXFHwskqCA2TB7YZ6/O
8hdilLM/IwhYte1T4cKKWA4F9S4FLrxrM0LYtMN9gXjChK0+C9+0AhbIrSanADXuhkyGIJ4EcamW
0/v5CMBjVf8/bEEzUWFjGkjIaHQ0UBPhd6JVt0sdpkFLTRq/F5pFbW63vPFNrK+1px87VdL+6h7n
cLx6Minbe+Txvg70KFyFOtZHUMjrGobukGk7B+mI8h9oC/xY8O0FEyaAwYwX53qY9pISV1CjiEHa
O9nQyy4+ZNSQFY5neTCv2OZc2s8+SlZLBl0h5OJpKtwRBnI8sAZG4ZwQKrF56UA9Z/Btbg+g3PYK
ZEXVovR2HY+D1uUtFpjzdUIDqrCS2T7ezCk6IDOAe7jnmUe7S0IFgEKuTE7MI7mm1mICM6yzRIWS
PiFHM0EumSRXPJyszMr0sv6CeV7yAE/SvwlzM/jpk8MRzYxMOh4qLBUWK3IXTpbKL7SzbdljhI8j
Zn5v7qmlp+We/aL8uNztA6pUVVQSn7yhgWA99eEFD8CzFqIw9Wai56+OdHn+FraFPcdXffkDFzP9
CizV+pVuNuuxyVGi0R7MEL5SgaDoDvdZUZqWhuBHSD4h5o6m26OSr71+MoOcZjuVD5MFUuM7GpSM
XfGNpY/tX0b9rjTrCkd884IPjo+V15Gs0y0oRWE/xHqH1H6mjmj86uPPUDkt68dQA2DGNCBJIfeQ
RFR1l/eDZ0AuOPr1tHf+cLMFq4JWscDKahmp9uo+Y/8YVExjoq1HCRQpvUC/VQKuBlSiBtDbFsHB
ax5lmvP84cOAbbF37Ge6vO6xj3/ySk4CvtTrkDli33xaBVqKShST3vqy6Jl9LI9Zd16Jbozz5kTo
yUeJuw4AyNIq2WiOLDyUdwjUtimFe5WYyiqgu0B0N8WqUwTvbSYAcXpN2gHfHSV6SgkErN4HEuCg
uw8Xg5sA6V3lM2ii2O3Oajw+tWSpPlMMZdCZAJSSaL8qLss5T0gUREE7S3tFPjs6RivlUBJqPp+1
symMJzt2pFbWJBjKQQfAcBgWls71L+uOeB03yNFLLcm5UczZRvfXhXfcc7yzzYnMkU955aF1CCH5
5W1W8lpwGVE2IGsjRbxgtD4I9sthI4fiJnjtR9zRgNWqKs03mtNUOl8OzK/Y8M9KsQLiVEpUlX2E
9TLlu1am9S+1LLFnMfpL3wnalNUr6nXSvKxiT+2Xl0H7m1J9Vgyf1i+m9+BK73zcqpGh1X42ZUBs
ghEUrHc8J+7ycBQOhd+ActNeWcyxP3jbAx1rrS3DhiksOTjZncuU/hG2KiPbijuZgQCrrztSnMhC
XPtiyJjp94ndmlRtoTgaKdJpTC5Fe1B139PJvSqDe4DuKS0a+BWDKamDvVR4/qtHFpI2mfy5Buin
chJoX/346xDUzwHjZCT4sX72U7PYu/2/3rD7aSFi+MGweIn5oPx6jSdPjy44+/kJTaxXf+UhF2Zp
5VU2c/y1qrlgY3K8F6xRvJkkvkHSSlpz1baFwlIPQFEgyFMUls90NIwzZc/XEc9Q5T1fKBK+lvvY
VLB713LxQUhXWJqPUEOrfGZ1CGtnPseKtpoHzE1vNdMS6/E7ZKDZc4OBql20/RPIs7OkgdNZfjtN
sbJ5sx1GOsJ75sgI4KIvwcnsMloXgub63bmelgVc4sm8U+Y9qOrH0EUXbxoQZnGAYl5reWWcDbfK
cwxCUdnWRD6TKTc0H5AiYiF/rxHlHQFi8keuf2PByZeVDEw2BisRKtWcGjGYJzBEmRIrns1SuHd5
/mNmsJya+2nuPc1n7/sav8aIdi9z+1ZAT7Ku/Rbr+4caT5d33qYRC2hmMG96dWhRVB4OVuEDTQRX
RYvT0Rgi33617yUQu/9iNSBXlVpDY6sdpxVaxoOaiizACgk6sidRbu9z2SeiEHzCdBCHMnsI1Gen
C9XiBsjR4U/snVtyOu8+lwFFme4kl7YNsiSfR0iSBVC7FgKBNFry1hFVLxNGm7JWvQxDvwC+hivz
s1eovT9xFU2CzPm1SD36F6XXBte2bJy7kwaBoGwal7qud3f1BGGsHvxspWGoEcG/AWwPsYmmJk55
VjopIYXP9uCMmtutvxhdbNqPcINEXH/CfA98jKmfRKD1DTCwIBvlSZLY9dbLRv5IGhfZRm8AjKJN
q9OsnJxKYSN63sQgh5ZaQpZQvy3k7HEP2rySzZOZo+Z6jXVXiSNYen51OxXkn0zy7V3vxT21gd3x
UT8+ljkrSrEy2XSujpaq2jGoFb8tmkdLOA1+k3Yr14ptI3b264MStIRZ95KB0Bzv1ZsnpZV4ofrc
2y4L7HfuzxUAvI0SNlcoxmFYmpP5nvjX59YN2cqhmQDiDUwr9qR9JvkqqMWCarvVrG8RRikHzFS/
KFWfrGGLvkxL8Qt97wF5aTfXgBWjTvzd+nBI+BkbmKUsPybJponWJS/sApehaKpq6SBxLszEMlTP
xcxWdXO4lwPHGhzuL+5hxvsrlRvOlHXiziyOW7xsjaC4lliu/7F5D5x2cIF8TfwXIH6GZkNnF4wK
zq+9g0rvO73fYQR4Wami5IoGgK7mDDVjg9nrmPkTHerx7fBR3gdc6ia9EznjMzerbLUKgP6nVDkK
zAwMDTCh6Rn4y2aOrny36DbEeV4dF9/VJzQQwgJLYeAbC1ZP25jjnEqS2hhh8AMGT9/1KUjkff9/
2iMIhqxDoTAWgqwechJ/oLrNq8AQi0JoTfB8/+APqg4NxG68prvURiBEIgZp7RZJ48mZzCiy/G7l
/NAb/h4EXF4zNHZD7KXnruCpLA+Q1UtynvcvwwBEmsTm5PG028R6H5Q/xIKeO0pp1AL1K610ftJo
DF50PXjWvP/uzrKtWkuFWvxSmU6hJnsQd4JmWdMgcyCBCJT965j0r+8CY5cFeus4ZfptrZbOlDI8
d8eN6rVA3GBvWMx9NkG2shYG+Az3AMfi/wAe6jr0i2/ngEnmz94WFhsxfz2I39p2ARiiwFa9Lcoz
8JKQWIwLE6/Kyh1q3C+eSXoSqT0WDGFOlInHq97YAhanlHxcXmnYKv/gvvSwRBp3YeL0kSTdoA43
m2ycgnIPXKAX0ZTot+vktWPdVBI4ReYRHkWQ705SNQ4TgDw4uHS0oVL3e+jDPsnkeTAniVcw1day
2CaXqcbwrM5vjWXmwWqQ2/eTSQ7uM8hroarYYkLnPcH+98a8mxmZHwKKGi4aa6dF9jo1P2qeiYwq
dbw0aTY/rPfd+WESz1+sypP0uCZkFZuKtlP1/RoMnvtb+rqX2ulhAZMbUhoNfYvJn4WVA1tL/S95
wae/gL+280dB8tS5FtE32QuvMlunEb/sFTg1PM228gn4C3rZkcIDNhYTc15wakhbym20lOx1sjP2
tRHTu+aolugjPqKNbeg9eo+zUTIvk+IMq7+Y2XicHD2I9HXBaq2iYpFZZlgSPi1cMXDx+SF9/CY7
+MZDl4gEkyzQsqrK9+9pRensngX9aa6JBfdDgCnwwX388dYYeyK7aAabqDcIyOjV2oh34puYJsAn
eOi1tEkStNF46r8SDh9dhwLnOduaLHYrNF6cLP2HL8y5SxYjYnHkyGhWmmY4wIEOVX6DafsqreOr
rqNC+1yxFPOGdzaAiRqN4LJjUZCNbHQo9NunXjMXJfe1njYCMg4taWoBuxRLyRS1zdPEmQ00VdJw
N1HzdQq6C15J3gr9L0+M1Q8ifwlsisRB0UtgbaCteTpiaYVmuU+6xXJqvsxS6puJtEFubrI9bfnq
jAPZR/8LeK815tlOHv2yv860naWEQdh8tn1uhPIlywmXA5cO2nvwFFsIMzSkGOqkLuGoBahXbCur
r57a8WgPGlzbDqRF+NhY5Dm0CaIRb1mPNTIrQJLVq86JRr4YVH/iOE52y8OeDghWrn+3xDbNmJvA
7VUEwVzf9Z6nlOBl1K+GFBAHi3u0OLgpH7Vf1ou4QNm9UylPkvgtuURPd4X18oFWhQpI5Z2zSklz
pz9mL98RDuIvM1XoV9uup21KA/Dg9a8teIoEClo9DgJoX0BC+KTERdhJep/A2BBBtzNp78UN/+Cd
u34uNNEVg99fSJGwiHAm0W9TPOgzYXUSbIIEXI/8jDcxlpd+5pu4NuUfT8fPASUTvbJKO3PYY//9
e7CXJMpTeQROduO7xDB7pfgl1l1uMQNo6G4n4R5YUmRIO3+PRZ3aXitZgXLivwdK6V7UP77Qln67
RA99xPoITpk/mejarau/oY2I8M0CsJ7iQCFhznzr7KUWGzMOjDjGHbAYycW4a9hAVw7OeMmrBXI/
9x5sAbyZ4qkbeaC3ajJJvDC4DkZ/ozKTJ6kdIQ8NrXkX+M15AqPZw3urRZLTotSJqZ+rT3glHf5V
ChhRQHreNd3TQWOuD62YSv/SDuHLDOQSqlQQOcvlWmaPo7NZkw7Z3BcGPV+1va2iT9rd8xRiwJGO
ourjvLpjUk35A0AiHrPjfwoIgbUMho30hLCggtywdprDxeeVyKl0mVPKnicKDzZWBiUJDkA9hIk8
yyP3TcXvuyTJiWvKAWIpUGy73ZOaYcCZYwRWwPTC8kn8/emp4Kc1l1ms7/cyO2u9QsbnYApfk0h2
bKTFpG+BB2Rn/wecIcWj1Ft50vALA1tGckOQdwKa87gGeHqMK8ivZbNQcmpsZAJtlu/LOXbp8+4u
HFUiG0rZB9En2Ea39AInk2wyJYrDxUMfGDmeIF5XexCONG8guGKHrPmTuRA3ggRvyiUC85SI3Dhx
xKZMwmG8izQKD50XNxSMiVU7Q45X0iFtJFkg+CU7QhLH99pOeI2AE6tq/BWgNDt2SagDbVh8fADU
MK4j99xdfDDhBanRC1THyEJJC+Y64qNBjkirpysNKSq7zo3Z9Qx3La9th/KtHBh9E9or7SqsHnuP
iTPfZI21CU0I1eu6uEuH1zPcAX5fgKbqDQmJiEclN6nBEBuG1KzF7ejD25a1H+rglmDSmNIYZPv3
M/mHHc3/dkx+OfaBtZQ7Vo6CBfvEikGTgfA8Pnnxgv0Pel6UFI6MxHTvChv6Vuaqy/bSjeQ4CeAX
u3xLAjsSL7ZczBalQm5uWIpRum1YO/G8mFgDyLPA5jRk+PPw7M4WD2d4Ve9DEuR6TXa1ujiK39rl
Y3CtFMZJyu7VTW7PxHzLEOuxt2EWmQDNSFeiPQ69FR8l8LJHBx7uYYXc7md3kw3a2ynbAtSs7krp
fGGFaoQgTvq+DUpm5oRn1dw6mOg7gpda5CqnUUx4kpcKgDeqnY4JNJimFVfoOBDf4yWfSuHI2A90
ptZE0QjZlyywoLbZ4/FdBo5KlnM9INJLPMkDn9Tj30j4hbbnuNheiPGkMOCyTcqczhdLENw8l6RR
9C2krYnykL0maN86fSCuL15egczTrEGW4Fcv691tpBlPKvBBUOPEiyZtMPN7vhydK3I1IsD/la2L
bv5ephdjhy2Buw9KwguqTZhRZb2jBtSE4zYP27ClgzQNkghrGrp8iVE3CxPpETvpHoKu8I6C+XgQ
aUWcRs+USq11Hx1THrtpF2OSefCnghQZipdrOGiY5ACjj2i0BRDFnl8qkZuP5iBZ83dJIRhDtz69
igc6FKfJMrKPWXa3PyzqmOFwXrqRnuc9GCnysTaWBOOYztlU9g86i3fgiBvZdZLpSZBV1yXDZgdH
tpsIbjf+Ak43CVF9mrTFPYxGwhFpqtww5glwBZ5CuX4rwpl89C+woPqxYUIYpE4ysA9d41zQkhHB
hmuXEFW8qfFiDE5d8EIcEvMaOmGsCU8TfolcnS4JAwsGggssUEeZHFXonYDu6BT+jbH9Ca15fe6z
ap1HQMXhNafFji9mETE+ehIkL9BnjoDo+3VaPuqceu4PgXDD6h54PbCLdI/uO/mWVOr5J3oXdKWC
gbThZ2PBu3cFuMLGKe1QJlPm78WsVGcmTbFAOn8qI091PCatK5BN1GcbIDYBsPypCyIq8mR+q9ap
0mLoOM3D1o+C3kNS0gV9GXZZ881WnQGHKYZ9nIon31RoGrLYOBtgQW5yMm14dIXMcCpblisYYhoR
fGM33tURhihESJkJFDftPtjyWP8hBVaIr/vdtIpCXt3sFVxHMx1XantVnnHUrQ0E3n1v/SR1w0GT
QR11NomttkPiBQIlbG8Pb6DTERiZdW6iZv3sWXrAmXWeBFAHW/UNw9rRcSeKATmSrxBpzE9GZH4h
HGiSpwtKvqfg7eILq7RLXq95mApk1BkLGR8GmrGlgN8zM++zBZxm3yB4DI4qhHYG2/ihfLaIYTut
xn3pYSSHocB47zl3SMEuBwBDVGz2gV1XOXcsDdNqAsVCLBqGDH8Lhf61PtL/+esSTscJJgI/BveF
d3ubl/M8RwfH/iQYj2EazYKi/1a9+zM7M9WdKzteIKakMWXOa4IodNhCGdZ+lkpTwpWsCwQ7d73v
37RITh9ltCo/M9GuiiusgdSsqSgCtVWP3JUyvtjR9DRc+k6mls9MviKu8GDprcHPyL/pz25vfYws
43SlrfBtU8uKCpO0FKzHhp56I76GDETEQqBGOanlXlJecaeMo0ZHvN9R/fQW0uLmOT1MOhYJd+Gt
Ul9H4A2MzsVpbE0NV/TsylyeMbMZbWLbuunyf+lB6u2FBB4+dxPR2BGbklbkWL0HRH44bsHCMr49
mi4rkua1bwpJsmZk2R099G+Nk4DwGJRlm+d3KizZilv6iL+WZ3gXRsdUAnb++CRNpYdhNlUxEHxj
n/0KhZHO33dykUZuuHuhMCUZaz5ZiKLXIJrar2BQLWE3o+Y2KZkC3PBEQ6M0m1jkw7IdBFZ302NK
Wg2MQt3Z5UgpsmQ9tNtTCF45C3UCEl/FXSF4mJoSj3YPP8rCQ192pL4olkYtYnUBRh7aPRnCUVlp
RTwQSpUBDJBj1kNUS0KhD/Dym1BAdcsyRmztyc52JOarhWqQXrAaKlXbjjoygSgw0l8eAsEENcP2
xroKBS3JaRb9SDsOYsZuacbyHEEVdST98GKZ5klHWDB+2/I3OjnT1Al6PGiD90GLuTADbxMngmG3
XWmh+enZUttelAv5QyYGHBQ17DhzOU7sfLuxt2phn/tw94857xOBOhk5L9h8V/ikENv0vSPXFlZg
JCC9DTnKoXIF5ctJdJQ5M/VqR01hI60f4MH6UjKyiVvmfTp5WUEjuTQgzFTFZv2HOlQYoYSyQ2eT
TTkDxcaohdszPmSekx/mMNn8qgf+cWAhZeylH7cYa+Bmi/5sOvXDIyQRq5Vyhdn4jnBoxnqHTTvV
EULBt1ZfJHoj3anzzLyC2Ggir22s5pycr2a+vp5c7YMTCIG3RtV/0WMfr8urxkrlNLgl9qLhyDcX
eSKBuMbbpt9zGMR9JHDy/8uCqAaWp9SAeY/S/yd9IROrB6ErPsKR3zuxjlxeQA15XXtPvfECgwDt
QExzXkuX6XcWcEUyHsI6nKOt7bb5tH9CgZCf0hhkktvPocSMTXbOiuRiydFNnH4+kC2X8JSpO2TK
4waLB0MWxf7VeoH0xtwCfXS2OjyxddziBQ/8ta7tbEEu9n3ys9Env5d1oMjf4+yhsrUgJFDOPYSW
bTAaJfME4WTkwnFTtlQ5yPEgiHisHca5160plnq1tJzY3Ry1kekovj8Vld9DPrAtBxJOgveoMwm0
8kOS7UolXS8S1xk/GJcVbLUe7JXaks822bACrSP9uI9HnUytq1K4LgJmgwr56qpAeihR0132eSON
QbK9xooXBqjuiwAraVpSBl8X4jC827Eoet6GKrkNqJ+0HBwNN/bFYm/Q+oyh1mcme6DOSzTlZoxA
x8QPUlrsSSkr+jXBei9+eOMBa5U+xZoHePByEg5LzqNypRDI1hWI1Vm98yaCmu5w4QFt52bSPIWe
XHYfJPD6soR1s8X6D8ox8wAOkPezBAUrAva4IVQsXTpwjkWd/RUf0fnq/35kuYy0f25siCZOfCTd
ceKQg4FRk9D1LfuKtumkiF2IJBxkmtMddB2T/R2H1bvoBOWxrk4r4ykkdM862LDhk/Ds5Z8CHaxL
IYvg9NnJaNFSFeuQkXXpbt/jprwLQ9bYKOA5FBIyFuRYfjSnvVeEWp8E/0XitSa3n/UTRxbwEHfl
HCLXnqQZ/JCRYilhoEeJToAhSdgFWBcKdNKC0q5cB1Zmc6nSDdNHoqZIaZaQWgzozQnItoVfMZQm
mAy1lcI4zEzi+xXQwHj1LNbCzP5BtoZp8XNnWYTxJvknzcju8sl2I/kOrV2bFx4q/dsK6F0dYh14
R0lgVJGCKhj8KqMlrZCYxC3JFU0ZCjSWYEbzUi9E3f+S1+r2GxIlHHKygYDCH7uRlkqf9DZaPF/w
9A4Qvi0k/15NXXphMLxlUzedkscviBINjLLlzDr0nejMb3bot1lQZvxkZmtIEnt3bxjInMzZpgRB
OuoRCDTCxqMoEx+g4Irz+QejBLc2YamLcxaED0PMUQibhSrE6OQdHyy81B8vs2zwOFpG6AZGocrw
74rbOijwLR6Dl/VAzLhNRNBnXpybS+AQlRU+de0+134T59G1i6MVAfbP4sO/mdQiy0gFdu0MYzkD
n1P08fx25OoPbPeTwLofxgM0drT7p0uGJETKV4bG1r0s0uZGMfSjr5NO/bGP0yu8lFTRH/eR9TIi
J0Jaq8/9On0JyRlH4b2TJb3fHdFKjxfv31YMsqy9+7ZLGFBslKr6ex4EJj8UvIqtYsRAA6EHH+Y5
5/tJi5F3CoZ5z8llixBMJbgwb9k3qN3XcSSyvzfsVn62OvOt4E/L6rYak/vREiUbzmq99HUdAv3y
wl8F/bVeIHJZFguc7g==
`protect end_protected
