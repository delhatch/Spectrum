��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^Ewgh~>Q ���J�Z��Rt�����qe�Ғ��/�^�I�	��)�(XUi����lFQu�U���q���JdB���,?매)\��G���b�ua�G�:����>Zx��#+�`�W��x��[���Om���^_ִ��8����0 gUk	�Ue���n�8�)�8�'�O�jd��AȪ!4���I�T�)sb�|���+2���J�5�@���:�� _�a��!���jbe�o� 7��m�=���̧q����:�y�t�9D�ӾVr��ڍݙc��z��LzS���v�s�5u�G���4җ:�����Y�A�����J �3׈��v��ʇ��suXf��]�Cୱ�6go3%�lظ�?�|�}\�I4&��W�!Z������sX��6���g��B����覿2��Iʙoy����
�p};��)O�x�Im���2B�Ȍ��G����;>%`����*��\�aR?�Ɠt���>��K�2g�lp��)���{�`d�O��e@����L.�4�,���x{� j���䪤ّڿ�>���7�ȕY�錭#�a΃D���u~6夔�m���T�����u�7�ؕ��n��B�ި����\���>e<z�"�~Y�w ����8( juw �T�����"��4=��?�U.Y���6��t�Ô��t����2G���;��=]��mc��.�?�\�r�!�.�'�[�j0?�L��n�h�slϬh-��F�C#zI:0���7�j�m�f.����M�+�l*R���:bQ,��M����b���Jm�(H�Ϲ�`�Zq-l>����³�dLGO����&9���0F�Ȫҿ���6y2�۾����X�}�$�R���-�.����������aC���};W�D�*inZ�q �UH��0�����sK4T<79�E�7�=���8L��*K��Qn�w�u��}9��]ٽ���̝���,�	4��d�S�14�C9�k	�r�.����mɽ��T�����@���a��W���q�@�10:`4� /ܞ��e��R
2�o|-���Al�`�<M	�BR�4/�m͗Z}|��(2z��#�y�8NY"J���=�Br�dÝ"�hnOH"�0l�B4��0��M��{�e�³O~w��m�5�J��P��&f'5(��.w�b	`�������泓h�D:�O�.y�S���y��^�����,^ r��C`�! MV�$K�kkn
�M�D�mj��?]襲����*Y9�NJo�v��<��9�:���h,��mW��`���?t�Uw㖷�#~܄�A&���/i�2u_3�|��fZ��Ȇ���8#6hx\�ﾊ=C�O2�TxpV���4���]�g�6�g�uh;>{����h_��Q��ێ>%�Ōk(mA�R��1�8 ���4Ky7�{���;!4�
%�T�4�r��jL�/w�?�H5�|���97�Y��|w��x=ԟ��Ǵ��%���`jm�7܉�UB�����+�s�r|Q�.���vƏg0��|��gey���1��&VM���,����?����tc�=��>R�|��uhT�^�y�CJ'��h�.З��T�,L
6o��mV�4�L����#6�~�P����E9=֨��RNɡ�)]���=q��_ۉ;�S�/=.����D�J5Fl}k4��w�L�&��>���Wm]���?�$4���Wa,��T�wdh1�v�uF�써��Sh<2�Kx,c*v�w�;�}P�🭞i�ʷ���=�>��Mؔ(RoXO�<��x�?6a��������a����郕.�̦�У�
���h���|,�X��,��I�x�1P߂0,���_���h_z�m�Ʉ��ǈdE�Tx���k����ax��ʫ+07咀�S�0j��m��ऴ֕�4�Ŷ�^ fj҃[͡�,����(MzE�*�r�����No
%d$a�(/Z�f�ؑll�G��x���D�m��	TT4�꜖�K���h�!�݋S���VQS^��:� �;�m�BJ��>��QQ���@����*'x���S���E�3�s����w� �s�X��%�6���/����дA��7B�r�H_16쏼�߉o�j0oDD�@tJ�?���A�-���;8�d'݄{�O�u�V�(�3>>��N�u���.�