-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
N/KGrSoF6Cq0vPkFKRH36m7Ih1Qh+2Rxu4WihKph255RPTbq+foTFChdsx2Pryw9YC6c5WRN67+8
gV/egXPGyVKIGZJ6qRi+56wQ5gmAQvVBPqEm/0W0Z2r9ki2acNG/CbT6RDKNznLXwVjrWUPvrVX/
VDMl3VLcgHKDT72Kz/mSvC3AVjwgR9wIyJXo34506AX9/dGau3WnuEQgDcp39VoQACu7U/dHDO/n
PlMjEh49j9zJP3AE9k0ZJv4A5XcQg4MU7OAjesXaLR1EFhbEZs1g4bJKMNIqhHjb5o3IFwCl9o72
fEdwJpv66nxOiWI5ktfImW6VFx6PzXahR+4Buw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
yvO/jTYS0gz02b7oQRkpvFK4CSGYUNsDoc2NdbtKds7ESbWjCzgYM8+WrSVQWiRyCNtD1aL48p1v
CYmPXPk/8kR8Y01eMO1i/4Sw7+QSRDbQAdQ/zI9ptDtFINm1vx1CiQKo7AIWtqDn96ALTNw06Qir
JKjBsfzNi1zwqu93LmhePq7HMKXPhj93EpzimYAokeJ4XNt03gzDGHt2HepK8L8298590hZgLklg
MVwUpoQYXVFfjC+w4GmaqE1+7Q2hni3Zffw7GL3TS4pD1LeibsUDXY/qiJyplIyYZn4U7AU/4oZb
/DtwiIIqzA2yJoqsa78RTZ9fLfRsa5xrHkA/aKrpCcgAdA7b8y5vW119cgp11xF+UcmkmEZblg0+
qoZIK2oH+fQzphINkWlc3x+AHseU/H8sl4t4ebmNzzZytCzh7j6JCtFsRRlULL8J5VygqDXyMZgQ
ltHOpA5gWOSh+rIBqJVek2jbX3S7ZIX6vzqHmtFpclUzzix4000QiK1NLGRikZlAY3ZciGXBFiHq
jn4OyqyzznygWRHaSaE7YkFkTI5GIyGtm+iFGuGt9cY/FisnU4+FdtqZlHruCQ8Kf0wBgFPj1DAI
YkS54eV+v7qh/prLd5jndFxZKr22mV28fcz3+lhR2Sjz0L1iIUqSbQQOwj25ZANJXojCo09YQHwZ
ArPXkJWbRBw8JBXDV6Fq9PkWqlw2EnlKmx1ilv39hhNXbeJuAXJNaSKtf3VXT2Nlk4bPDWirGMYk
aJRg9Yx0JjBMb7FVR/GR1TdH2umGm5mWnlEtRFal+8T/V/3g6oXdfncDDolq3VnuXaqkJGTMnITt
hUD8/7aDOE13N5SuXRSBabAc6wJonG2CrywsV7Y5y6Nnq0CL8Ef8GaktkkHoUZczOuYx5KFu+LF/
9ZYoVcn//OTA3M5BwDvhxHo0Ubr3XeQZLtVWLJ/lI+Q7wQ65pYqdJYYORK9zJ/NZq6C097V+Qqu3
s5Q4fiGi8Vr7+ylTA5IRjFNmPq7I6avE7L8/xAhDnSvYI0d0unBO9pmO6Tma3uczH3xWkCX6WDTQ
FtbJtGUJMVFqMEoLcjgMO1K+UXKUbD1d/Oysg9dtw4z6cGpjtWlyHD5PArE6pJ2Ac7BU/qzcREkv
XAxuw5gYeqx1W43dgqfnFCnienY1s/mdrqFL7v/6GmyFPEkceUUGT8bR2BgD2YF4MXxFXHwhdaiz
LsqlmLicHxaE17RyCdDmxVtZJ5AmbH+7RJEiwYKdr25LU4psy1ZKAcxDgA+oaQs6w6nLxTro/G+v
mPAUjjuBA5sxQoOsl5E7jUi01Vuf2Pi9d3U2dqIvZWt2VqLv8pKG5Cir87wOVlIcCQ6ynW2ADH4o
jVKAD+SVdv5Br7fzyP+Yz7Q+VMroUJJuTLEEDhl8ZtSS/cI+dxQN+brJEJ6ZO3+dQbWQPD+rfGFR
L7V/mb0mWxhIRlh5KH8LewrVamkBXAUkMddSkdiDxcXp8+A9qqRH06uxNO43AKEomDXTeLcGrpeW
nB3BWr+p+Xy3kZZsujUU22Qz9mh9S8iCvO4lzdkP8r08+naH/SvMurUNCnGbipZVo9S+RuUF27Xu
QSfllXnhGyYWqiu7M4SZIYF0iZU1V0nluPl1uwpowCqdQlMgOaqurVnK6CYWXTlZSlI2m4V+jVcW
kui58w4fu04MeespxnDYUMeyeowhSntGOmIy3myMKqhsNTmB0AnaK+nbWgzsh6OFn/LMhRERavzT
8EM3NT0kvGnLrbISxpgF5vZPv9M27jmgvqyKs6GEWPqIMfW0ZBVXb17O13/eC/5QhDGQncK+9omp
IgmmjtNaNhAAiPLU+Ji2wouuxjOmEBHcp+QV65NeFCLuM8yX5fmSQ//0Lvay2dKTyzyjfjoPQx0p
LjEmXeetWoDxcLB2C/8K5cqG7tCTeIKeIHOgaF39AnjJfJOJWrIYJOadJRwae9lJkTES8Bv6JvK8
YOAWx2ebA/pnDhlpgfvahuKCiYm8UpK/Vefzll1u+V8hbeH519a5JpgqYylijEJw98IgUIkIALe3
fuj+HZ+BFTqTIoGpmBsAMWzVvO955j91MDknGF6Ezme3XM8KLkdGENn5tUss1JmdXAwFplLYCCLZ
4/scZptBAu/aA9m6aSvSNg1+5xdH8MspBEigyl+l/AD21ZkSxKxt+zDpTfgdf5hEx5EFvZGgAmAr
L9yQXADTMksqiRZHNvpoa3CPEWCawDpxed/utWBOsW1bDMccTMQ5qc+LI/b8g4aiOeXMsM3Ih9+j
JiLhl0rPZZrRxn82K8D6o7R3lPBBbULteNdq3ckxjGK5ufXc8c+bjQBeaBywgjnGDy7VFZyhkVwt
meusDaPIIMpPCvEfwmpblJ07PyLwLXFJchNg53HgpvWJZMjBy/zMmJKx7vyBttEq4WPeF0BebS5M
cb2/uoa50qFwbiFxyhVb+8awt7uMnAtB9l0qgro21TOJ0sl2sdYjdVveJE2s4ywkHOBqVgBgz/oB
1s/l79+wgttF0HaDeogfcP2QioDYC89nadSH9kKLc6SI2leWQXS9LvioMXmQmo9B05WQuvIFvDua
ChN1HrhZHZzn+vdgJxxJQkNq2laeIjkVlHaijcp/wL/vZoD/SGJvn4Ps3R5zboOogl3poTNnqAgu
V+JbVy1nTh0i8awgypfSjLX1tsaAgdgtRbzl1tT4Fdjs41q3+1n8h/vmg9BclGjBMkGJe9ngRUlj
CVkFAJYMhFjBabJig6uB8pbDL4bYt/Zb0uihVcXrrbKZ9j4q6wC1q/nop77ihggoTtdGJ39u134v
fzUOPuPXEtcBkE+7hwYqGZrt9bOBZDScZ32+7FtCsoCQJM+MQ0EUAaZMOZhsh6Wpd0px3B4J4Tyx
fgneN9xPt600rXMMZTyfjNrHKYUsAPVeg7Qez5hrIYwQ1HvnJ/FOTfjc/2CVfiSbVMQiTz0iR3c3
OGrJRbWPdjz+C7v4FjU+2uAgP3JebBjJ2jGkCGIbI8lvHegzhowVXVAoeWWc7+VQyQgIOA0wufgf
+pHNLBrN3IcmcxkhtosIk/8khLsDPbaBQ2njYbQ09yLF6RILLHsbtt0MTAYUXhJLWlPNFjLgkClo
BL29leVnFWsVlim4dLg0wpTC7bZB1E+4sh9XoxcEr+7UkokMTawg+I9ESSlYXIKtlK5v1nU9OeLp
1OwlxPq/9Ua1UWVPJnYWZMbfxo3060ZCPhUEW/1hQZ27bKfKktv1c3qs8raIF8+ki/8Nb4Q/iKvF
Lp6HDBBWQ2cnL/drFRfBCu/kPGOgDXnnRHIVO4cOoJfW7AEU0eGS1hvh3V7HDuzzE8LYfyWCZSfP
ONSashmjV7XnbCqQ2Ufz38v4uscsCUD+SOLCwv6CBJULVsOiLbDo+9wk/9HDpggGDuVDtc/vroe8
9Nyw/5w2uAIsBRYbhz8clq+VV6fJUXNA3dCl9vdLESoE18CANsoZPqD2x0wQ6CA24S6Ro/ubbQlj
s0hbV4kuH7GDwNgaDYcJtWSJm6Kyr6rvE3lqcbMq58POuaAKArihfLlR1EfJZe/83CTHb6oBpOmi
cQ6anjCJ8ltEBoS/WusqGviGZsoEuMlY4UtTbKZjkb41da5iNhVWsevew7Zmik35DlLfalGLKFDD
aqifAM1hMgTw+DsvSac4s9kuIEEz8bVAhYYsBSeNxcL3fLo41qWDEPuonyi4wN61WqEV/4gaFWeT
qBdQDuCfVG9vjD43mEKa1S6+jhnv6Mx3T9jHgrpe7qZb/eubkEpYPy8P37TSY2mUKQ11+HTTeH/s
7Mwfi7r/dd6gg26dSOjlMzT1JncQa5DfTfN4D/ei30CaOjJldcQvozunutBjuYx+3uqZA/oKWSsw
rrht68o7pFuVXeMz3MCkKv/96vwFC4LeFTTZO9KKc6q7LdBsfCQBFJ5xxLQZ2sLwS9wbsZMl3dkW
uxvIcrdejiyW4jCeOlt6fAY2U7B3KpALl9g7VgZxKfiOgfxunqflGN8xMwHv1DgBNp6qZ50STvac
kSYUBQHBBoq98B7dcK7mCfmkxsbwHwJq7D9ry88Mu/o68qynWG6e8Uvd7C5XepySdLopWwlqLF/e
CBtmR5Sai9eOyvN/d066KUvnbGaE7VOsIBJabrMxQaHlmGL+C4fZfMaAkmzzmTy2+O1/UvEF3LSr
DW58anRAR7rLeh/14glfqrCYIGQfcdEb5k/D6NaAhdyRFN4E6Xpsw3euKFq4VI0RUp2nM9t4t3MH
7MxU9Ae38S+cZRUZCvbNbdDYLpXmQ84Ju/Zr5o5lEqA9GevoYDNhsqDHEHkfe7Ux98ukvCIT7YwZ
LsvXzpBPe/Ga2hdhq+VR6Nyb+KMF35nD22rC5c1AvIbj8wkJLIYQFoTAvVG/zLEWegPa25fgHIrl
bETsXgUG+UjDjP5jXY4EhqTxT2p0/CA0mCrkSaEFJJ31xj23+YNGO1STuXhG7qujNh/NvyOWOTUf
A8x7m51uETHkbYTXBeWYXsVH3M3a5m25n3bR2Vrb6Pgi/nzwdplpK/2J+D+4f/0FMG+cKiiVAAjX
ITUEor8l9KO4DOPX0TiG7c4q9WrIBS6lt65EhdJmMZsbaKsdjhgRh9Qpv2GoyySBiRBLf7SAouRV
vsGCBuo9JY36z5B6mim7oB9cwVyasq9swBR8Za9tIk5DzBlFcQIJPuSwXs5H6LBn2WoneMM0Ph+h
mRFT9j9TH5ETt9xFtIj7P8pWWu1jmNoKRqxCrelYFpAW8zv5xBPw8Er3WFzWYEW4Sd1ix++5vCT8
T50HM7HiSc+iq4cpI8eovQ2gIQiLpcvEqkSSz0o3+sKVXVDSbljmjwkV9ewhgeXgR7+jKQAxIVxx
q6QrSUppvqxIzNjRTjBK2SdYD4BbEWVd4ORY13NykbdJowGdpnWUD2WPwj9Tvuc7X/km23v/5hup
hBHK+amj0/lOcsLaNDOeRLfCLRqxZ5GIhvnxh/49QZhxlGdfUJFkiFsrVNGa1C/+HPY1RvA9kRju
Nl/mWBOv/Gf7k3NRq6aKLYA3d3ycyM1+0x57bBksUPCrhvfyROj5nHJV5IsIAekJTFuh3CRgOqHd
p8vu6UUARMQNMzxvTDUE+c08S7CuJBGHKFqVZ9kP0+MTlWpjJl8xlgv/iMX7FCJqyZBPmbo77/9v
0KutYLvDKUy4Y6xR9TsKSmalXz/GYNXZqIwrGICiJBN55RXDqCCsQILaSe/QGshhkq5QkEZNiOJk
DQtIQA8M0nSJYmHElbQT6NVSu3rllmYqedpepTc9uuaTtMGfSAfmQmVLFRCTrsurW2JsQMGEyq80
Ut4JH2X1f1u6M7zxei47PpLeAZyWUdQL/A+wTUjVrP3mk+Ps232N4wGARFErINWh6GkL/PZca8td
wqAl4obuQzCoJl0T6d8gB0R7ndF/D0g2zpv/HB5sTQeE3g1PwCA3y0DJlpfLoRuyNkjjBxg1efRi
Lyu3Z8dm5aBiKhy0d0/mJ842hi+0AVlyu0XmjfnD3WKnHD4np8E1GCbBv9QDKrlrQDFaVtDI89M8
StBc4PgpCncNdN7ymakISJs0L6d5r4fUGdU0uxQMKAsv7WqYI6LWbQqE9s/hg1x8zSXd5TD18CN/
atphO9qG1Ki3zHBSzqyxoqgnBWif4RC9EpBxgvV1w1nItyf7vYKZPCE7A5z5dJD/iH6Dx7MOXWNW
YIK78b8p4XZc0PLw4wNOIFTOVATtZ3a6Ivv+bPAnjtaIGOca53AnWX9wCBRMKllNAyGUnb24ZHmc
RiYvCC3kyCQPGNDXTGb3V848kYfSzqzm7WIndzm6iIywYPfG0YCMaL/rO/O4BLZQNDYPzuuT9zli
g70dwHtWEQsw2VnS7FIT1xQE3upaC2Tjv42L1UgpgIIM8U4aHD7tsKMKLTZ4Wl22I78qAp7wvAif
cD4KwhAailjijYL2bUWXaJ61mp0kpZdLD8DfG89UmoBLG2UVoKHp3DHArIAEEoxOR/16PViJb5LK
s56+M1cftHBHxcVPNZTN69ib2lfw2lBe3hWxbnhjYCP+m57zHuPJ4Bd4pd1K2sEZuFH/G1Btzb/H
1GxdADw36xH2fKaJPHLIoU+RW2ONzTuSulAsoRul6g6Kc3JC2eAzl4W7/QOAxVGH5yqOvnkSRgVh
WayinrXAB7YbPlBxy1FicQ/RNSCh3wjWeroRPPNBlVxYnOgNWx7ogO+LJDZoYBtIAaoA2AQtfd5t
Un6cFUGXa9ubuRXAOIt2P5oFUoQfyiPANX3iX+WvKBdJoMt8dU3vhuGXh1jiC43S8kmqJY4ZY0F6
WRl0dWUfLk8UnBZd6AwT3fI4cTyKxaNwfiE8uUEjw6/k45MldTBdxrSj448KpVBivdp1tkeH+jiO
lVNrJhSjUgRKEVXwxV45OLDLc3m32FQvSkbsL9MpAsgJv2iYC3pkLpr79cNH+cKYi3NoHiC/5Uid
UEfOohKmcset8IckV9X5wEMcIZx0EpikTyRBCXWvNT8aEQgdZDLVbeWzzSiFSkmOEmrKbnNSrP8l
+tQGprHqIehj3pQ+a3hKpApJgzWIUK+MX1LFag760tB6LDQVpyHJhYnkE3oGNCuUtEWAuBxhbGGd
RDBilTcwaIlc0SW3Zan42g2tbPbQ6BE48JAjtw6aUNKfNyZe1BIIHRV7CsMRDEYoxj9Woxkaixe/
F0r9y31RM65jZl/o4EZl4esseENRmC14HvDpRRt8foVR9edv3+WgXxToCER9QLwDhX+LUxmxqAGw
q9MovXSw57x23uzSiLBMRpBLu1h3aPvgFuYFzZQYSvXPG5zMEt7sa14U2oKUAatW2V3cg97JDYM0
BkFCy2K5qPYarhU1xmbuBQNfJ3TXtPFl8OB+FDG5YXZSrDYvSzTSo58HzLR6LDBlGpBxtnA7vRQa
L1g9VqNZ4lw4Wm6KjBTN5GXG12rrrigAYaSU2Xi2LZMh++8X7DByMhOof6wWyFOcwhs2gTIo3b9i
SdxWTt2AjA11VdcwU9BZ1XCerdw87IpscXdTQ7gcdaMjp+gYnps2RSOFw/DjA14lBzCEh/St+0aL
BidqknOqygh1kftVBhCJbaAnv3ZmFsSV5X94B1eKDaOLeq5iy/aZ16rDBCi6NwhsJQhin5NAH1wV
jDWGcrNXdXAu+xxuHi7YUWFFqFhXmiPbE1H7rn9PNrE2qLKP51kzvk7lxcf55UIRW6K9K76i+dUb
ob3lAp1z0kqjeEJwD6RgjJDoHC9kMmr5leD/NmvyQSFpfhr7kJfdNn7ufTORKOn8oVvtJUwRzERV
U7OxJWKo6In8BoBEVaqfA9YD1anV1gQmOlZZ2B5VTIXOmY7SGzTRdsewpm8P0g+B4ShgEB+02Tb4
Vso9KQnXLs0MPuKxU2YzFPv/yFF37hNY8GxZM7p10hKUFX8izmBKg3T5GpZtWjCjSDbuzs04WeBY
uVo3jydrU5e4HmDln5YTsCoqsIFMhJy8LxV8BQQFgJF6KfMbwzrzc5Q6KjB6OguXgfQZHyt9WYi9
xUxn0tsM2C7siGY6JijTL7YGTapcHqRKHJeaSdT3b26mTliU2pmAv/pAgIplQGkBUZ5hXcajEPtl
01fKzOr7GvAxutlvlT1QTjqh1CUOo2kRMt7wzjoQvLnWebgREXK6vo4IiPryvXCXX1OlYg9YGMCm
MRuWfwO30TXsEoNlt8M1bK0tSDyvpBZZRg0WamfSAjFzsl0TTWVDXq6WORlGCUZ8qjrrS1wJbT8m
+j9YgZF1bPeAyVcFTawAoQe3d1OWV7y3RSGo1JImdKf8V8kBrb+rAY/EauD34A6/sNAKSMPEdtV7
YJdw+5yhWhdCOIgceovQkH8/xitfFj3gZB3WyXYsxlOa1qBVjox4kjK5vMiMpQCpkArxxW5OU8CZ
PzLNa1jvMBh+ZgJQ3I1om4Ct5cx7FkkP42wHLKGHkFSDLMpbEDBBU6H5h+yRClERR0OcFyQ7Z/4D
vrXjXMzskWTXcWtMAvBucbPInaC2LCJssgeMcSkK7KtgBi+uT9HWR6JwdYixc86dLEgAGZvqyLbi
ZZ6uvcZz6az9E8OpTKxswR+qaV1AADqeJIwy7T/i/QuR3cdlFiO2KPpj8/lJvEf5JkqiAIthlBjs
SZkjvl4vrhYDHsKY80UJleSAAGMdtJRiz0iAZvSvAubgeIL3ZXB18vLQ1SwGmzH2gteEnCOMizFd
FIgWyELxulaBGyr9FZsPLgYgzzW0z3AHbN6ma4TJhC9orizxv8wHTzoLGLI+qJgfyTJsvPDSvzvU
kb8lur01roMEpw+E3FqVMtfUbOu34B/EnZhUPZaFtibNf7n08s84vD7+bPzdxzHgGAsyZ/oj+bxg
ffAkbZ2zbbWJSD3XiNOQS0XO2R0K3ZX/Ky8c4WI6m/ccvwu1csiwNkVfalRVe/Gqf0vQnuWeu7RZ
o5BOMRrKDXTm4G1voCxe1uA4IRF+BSHpl9Vhe3YZPY4Mu+Y/zCRMBtaAXg3nS6HJpDqSKHCFhrjD
Jaf6Z9Lzfc5ZX9Jh8q2BmdNtB21tCB6sr2Vzg+i+5x7DAURKZoR5fD+nZpfmMO7jb7XXswxRkJpp
JcQIF3yLwQ5/oLqxruy+5/TZV4lYKz6/Thg8PYcpsFv2hED0LdhWfyzRFpbZIvWl+vhs0grlzAdo
U19wLbc7GIXHIxehBJ41WkkR99de6XS1x4UqnepcM/+EbDYOcNkxgj08YY08/a4B+PiypnRkvWuo
C569P0goGpLoDNvvK5eF/j1xY/OC5mEYSI0K/3QkZ2JtzKnoRZgRBIyPobSCDpkms6KlR3tUYM2h
o3Fo4t3zPAS/vChtuiIHZBA3+Tgo3We3XU94E4pN1tHk9eMeTiG5Tsxdso1qpvHK3XmRQNchSe4k
vuOxtCZi2UQK7gjIQPgH8SA2rMoUsgSLFp+fRh37aMHBy/aVrIF7PhIu1WwNh0yvQN5t8HQ7jf9v
O/Ju3KgV70MjasHe3V5MMacTP2/fsA73pau+W5sQWGybNIRCe5H1YPtmr0IfaV+BQEHu2nCk4pZu
vryd7FT3AGLNQ89QNI4z5VwMJgSazlWvux77eMbmubPC5kPGeWvxUFT7+YLx3IMweoRRC2LjSGlz
w1byRRIbBKtfC0IAUtwK/Eeb5lAf5P5FxqpgOJrahNtuQveog7NUbXG5sIgo8hFxv3aNjqASjkLz
/+od2s17p+N+lMbaB5fjQHGSeRJrNXY8yvYxRggkTo4jFagq7bk4ZyS7swVuCU3jw/o3w6GtCEf3
de42t+u4eXlqFqW74h5672/KNJUAxqRI3O0qX1NwIEc990ABmosQG1vSpLZuDlYRCv+KEEKKtmAx
55Y8Zdrj9zKEO6aM7sXLRo6z/ToLYY2eoymsI6m/qxDagRrCzcY5CkD0l3K9WTRm8kHhVydoSYh+
NEiaQD1roF0EA5HvSzAHFsSfOeMdQ2u/ohV94wvOMEr0AdUUBo9T5WTzl+0P7RB9rv38QTM/FkLh
mNxpLYV1iJgd9VI7KTdXV9OiEkfE8LZcbBCZRg5YUewS6tH4/qYiRUGWqG/QPOFpCMS5Tb+tJoUA
IbB6scQ0Ya3BidSftcEJGQh6bNXGStGCpysC8it1tHk1aVK4oLRaHtarn8jquWlVW7f4CX764Bq4
RVM7Kwv7Qvpwl+UVJey+u5BUV5B4PJFL3/S2I0mJh7kEvsxTyD0PYmOCHP6LOcj9Ql+gRNQoS+tY
6eqYl9g3P+jKF+0NO9fI/cRBqLtNiW+H+uaUQBRTkT1RARFDCPLA/gZ7ltlzNhqfm+rPehWi5HA/
flhILbf/jGuOrREV9BYxCNR+C80165kG257YMaPURI9XnJhnbMVZNXcz66/gLDUXThJNSZymFfeB
OiY8loosCRvQhWbm7AUI7aWjYpK4vaqeykKUPU24h7X8V1WGBzy2uUtg+VREpw8SIb3UZcjozrxu
sJfHt6rfECx01qSE2Ync4BveuxjgkeCUS5rTiVH8xYOh3z0I/7qJhKD9UdxqZ4EjmSRnCXwN5g6R
LQhwsE39y7cmI8aKlIPYZztXf1DmJMlAnSLW5/dArQk0quY37zTGoA7vc85aQl8B0cC0/PZsCyN6
Z5kODukFn7egMTx30V9bRMYYI5t6In6WYDy5Qx612wyK9+tqxz4y9Z18A6oGlEHQy7OiSxhlhllm
Xl3kSDe1HuWO7gnTlGqQpxcgtbij5EWXgh3lkf+DIhjZwxF+rZ1gg+KQVmr41ksgEERNNmUFkQBN
4tJApqajVuzrzH72Lnh5sLYJkKl5U3FhvdHwzErCvgMZTt2/LZVa3wTDK+s5ySP2V9WHsiCT/TOw
zDQc+M+ktZyrquePcBAswNSAwkWPePHZp3qN+mRsgCq8v1N2j6zMN6n/SAHjVPvGMOQSt046Fi+x
aPU4rev6HN3gy001xC08wDaoFZURw0VS8Y2F3+1+uN68ug0NOLmj2S5tdg+m+UTlx6IWLRSUokUp
xPg7L8DuMBHnyGTTrGyH399ZT62n1mg/dXsAD7LEpAl4ZNKTDbD4PcuPoRXol9kFfdkxeIn6X+eJ
sInMrS8vHsrXHrY5pdyv4r76DuoO11XdzNQ4Mlr66dHxfKhxdMVpbKm1k7Yg2irShj6bfJrmQeih
ZN4WGi8T8+A83d/Z4J6RUhQFunrDQOVY3L4m0hRDCZmMZ/1gBVZ1MCqZo86Yio01sDAwGjdV70se
PPp0F034BmXVKJlnBzmz2LfClgyP92d5AMUg3vdy/E3JU99OUKUTwT23E6yRHkro7YK8qfnJRBA+
VX5NPNMMEZCtzrp5bcoTQjM0pK/Ipl2v3ddfOB0vOxbwZ866FIiJ45UCiMWj4xNgostqyDdMtYo+
I/nuZJxlCOqum0ansv6e/oYyA6TJ/xXWXE0ScUZOhOJpCdeotjfUX0UE+qFr6g4J5E2P40OiIEpz
jk+fS0ij8pQeBK2R6gjCubwvGUIYzSOjgxofjBjNS889EOCoZ1vIyeu1nHnvSDJJWab4WIPOkrfy
S91IXuxIcBu3oDltQ4g68YxiBAhLWID1epyAOl7ggkzp84Kj2h++LyPHMeOepPhTEm1jN2r5PMUE
Nxejyxh1y8WL/32udH0n6/h20vOYYTLZ0NGcQhs4DuQi/saVQXY04TON1049TK8JuJzT6Hp5fIwC
F990DFTGnbZ0d5EAG6kF2ISrvHDu+dI1iOMijtYdX2DAIiZIpLK8GD2Hs0tlEQdmvfF0wBMLiZLi
oQ+Hbgd1nWWPt+cZNi52ZxJRbVBlcVrFFj3rQic3rDFbv0xusE+FGJE/qRaS8dSYaJnqdy3Lo6OP
jT2Vqu1y/7NpVXPfrMj55zuxMasSo841iGY4K5XUcztb17rAHG2X4dg/XsBq3c2Wc3I77rUpG1lA
ADMZiIkCogv7+KaoWeyXTQj+7r4LoMDw3bcDcOfODMoEInfeYtW4NQXhj6hSpHJptyoi/bnmHCmI
f1mWiyCVdSLJxZM4ElgHVJY6JoYXN0g1rT0oOWd6wj2x2Qq4jD44aRwt8NaRnGe/KVRHkSOkhIJ1
3gA3SBdjikLBFxMBVXA5P69Jjh/qNhDaCD6xDGKilHWlcI1yCNDNfOOPIQMxoA11hRtR7A0Bm1zT
CRQFTIy3BFin0D09/CTzwRyUmDxmVnGF0MsXwJwKwt9FpanAts+0CWITwAYEoLGVwlP6ns5hQTAY
hWacghyr1T3oV6eRukwKc8uo0Y748XtJX8rnprwEjyfwtaRANxlQY6VqWNmGVIrIA/1ewifFHLg3
4h7fOx84ogrfEy+fuD1IeVUyJIi2nqwQ3DGbOb6bELklz6IlrI8D49o36K9hM4rRyqabcW9Z7x9Z
UpEZie0Afpv3pU/kreNVC/c3udeo5q+PlzeJktxVI2G0TeQ4Ta/bOamr00w0I8uNtp8cQLNIYG1O
F/bwv7ZPLWvLjBFBqpKqz+knTu/E+dr+uiU8RbmKAHqxsL2pVpPlDQps2whCqyjSmM9FEK7PHpYb
Snmrml42u9+DNMTvg5Lo8MjHmUE8FtPpT1nMzKvyXzfThQnNNctd1LxSfCwMP0GTHCD592fk/kY3
0fNpg5U9UiqC01oCdDU3zPmm5ZxjblkniWo7VMHYq6NsKFgfK2QSa0ZEm+/0gtR7jHMNmIYPMYF7
5BJLwroA26n1Pqb19u9Ga03nUYV+4E2c/ecUPX7IZsyRkArUZpJfat3IH+B0mx7GOT/MoLHf/KTA
rhXNy37LthuSegMtuk/2KMUJRdb7A8Le0j3u11yWeu3Q1W9c5RhNpdoiBD9jaD3Zgh61TWYxHrJI
mS4ISyVv+oJrCVHU+vydBjQzIkbXd1BaIlWN+ardewQy89LW8LqSlCvqHGd8pQNl9G67RQTiplKN
O9Hsqal0h+u1Q/u48nBHQ/D1wcS6YVWbEoziQa9yFgEWvKjJMr+Z6qCrfTNy/2j/W69ydW2tkSKb
oXxC6nBQq/yDWUN8jQ5JxwhRRg+X+/wWTePHsL6YOSX++nrYnq2lCHbyi+oN0B63rl8mywH2MtQm
/0sqHbXOY4+aNcZm4UJVZ53bNibVaIUoykz2TxGZ6uelVPzgwVRd2tKbg8HDWZL49zC9dzOeMhZj
c2nRj47uey/sAVA/RAGK8ndArpRr7xf9yQKAAO07MJ7AQPyGa8FTimDRpZd1cA4CPUHopD8wmjd9
U49+miJ0H72Khs9Wn9aALk7hY5sDr3GI7PbnBxH4OIa0oiPurqpGB2GC2zIGmhi5TTQgKb/wL9sf
GN/+LhQqIrxORHvlndYdlagrLaxsFNqUDa3yTti1xlIh+t8b3s30BDRKHSdbg+BMlTg9CWXYr0Rq
6nE47+jjF66iZGk7ArpeTMtAiJ+dktHUPSiVnOCBUK0Fzi2AmP1vkTEdHRSSkEpc+vt/eDF4+87r
pQSgMD9OHHbHkoIkrH11fKIb81GrICCcJZHu6dIpVpZc7MYrGkYPyh1pbi3QhwmESIFSMM9l988z
B84CNJybJ2lCzYFHp1krvkXmy0FkwgobsveE6kXyaGZLOXkEoNsMHOw4hH83/9vXnRsnKlJU9xXb
9EbyJ0e1xfNOaGzIQpCO5Ir5EBcKTqQq3628b/Sw9v839FAobg/T1nX4nGxUW9BpgdLyZJNfAkcz
0NPXDjSWBeur3Ju20JM3lFHJkljiMFbFF1C9bfi8iL+htrAAmT/DV0Nc6IByo4NH9RaZzQhJ47ag
qVYZmvR4JVC5mD/eSIPm6cL29jDA6EME/uOd6r8q0UBO2ZVA3KmtEh33CCnH4d0FzK8IDE2rjgRk
uLRF7/ekg5lNazsP416/CuvgqRSCIAWhhShuxnAsHHcDKelVZhn0AtWjAPNDvAJv0uRCxXsMTepB
+L42tudRco/HimoyZ0BewiQOvibdZ8ILxduytv+Wb+LdenjbG5Ckp8FEMYpK4CS/bGFXQnWXveRT
bpTsngLMgRy5ed1bmNaYBUEAHo4Cq0a4cYkgJIfaLrmlXNFcgtMl+5Gcjka/NPjR5OH9LeV6+n0j
rDzKgRU5VhFcOR3lMagEDoCN170ZsT/W0Z/2tcxipSsFA6LlKUUJU/ncnJa2By6rK7FCZC7PpUsZ
e1JBTLwdh3abHgIaK1gnq2zi9ez/BbwCyz8PeGmZA9Yq+gUbY7Dgy4J6tEPb8YP5Gi2OT/ur6ul3
8QsNCWSBr1kl5QUPS5Fr9hJvnLzfx2s9/G218+KFQpC69OzfhJoyTgzooBkmQrvNgtdAFAharCSf
GEpcRhzPo23MQ3/kGIYdlxZFRA==
`protect end_protected
