��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���'�ʞ�~|�A`�U���k�,�ܻ�zc����9z�n#�?Ff��w�Ϯ��^�����[�0�=3i̬�S��
5N���-)�[IN. �b5
��N��@<�"܄Q��X�q�E��?���^�Fǈ��������0�X���_B�v}����M�A���v��&�����r85�I�]�ޚ�Z��0�[(�ԉMr�	L����H�0{���͋�G &�.�ao�5�X�.��e��Bg�-�4aB��rCB�]4~]�z�q58}��4A�fr?�i'�ۤ�r����IٚK~�?�5<�� k/cM�׾�V�@S��ni�;���T�jhs��-;��b�Dʫ�3�$�'�Fn���A}~d�!ӛ���Q���:?Rl�<��*�Xe����~:f�+��*_=�h��)�V����<�`#Ւ���q�2����{i�\�dd!�ː����9�v��
�@��o�.ky��V��Gc��������F(�J�����������k������?gk����#4�F�0n��w���"���Dr���9!m�̀�q�7[+��ua�jy�ډ|��*�{ea�I�� ��]S��H,�>g����u��ȒcD`�� X5j�����ԄWa��U��]���O�4<�Zzr+$]o�ǧ�"M���-ZGv��8hR���=�8w��9��譆�?p��V�y��#��[ZK��ʣ��L3��8��X�'�)��p��quEF'ٟ�X�Kls��'l�����Yx�Z�!�*��k;tC�z�8��x�������U��Ie90^O�b���4�u�z_������ÐAVe�(4��%�ipU�O�I6����=w�j��;W{��xS�K��q<�pf���_��T��0�rz�l�I��b3h�"�0�EPqwR�pK>�,*#/��ƺ����
�dxg�">m��7����E����� ����.T�5��*;T����DAi��6te��G�zv�q���|�o�믕Ca�|�����ڟj¥=��ݒ��-HuO��/���������i<�N:#�8�S�w�{�x-u[Koy�FK�VwV���fŎb�F(�
���pP(�S��N�5��U��H%�6�ڻ��	�K0X��=��'��H��ger^�������U�  �n\F�%�魥�v�� �G���DJbMV0o_�|7�\*Z�v�Y�K)�����PL
^i��2�5�wL��>�#�p�qɖ"�7�NLs�.{��x���+q�牤�n��4�	[W�ר�|a��"ɋ^`R�S�'�0���L���n�δ����|d��o���x0�"���ތ�"޳�E��`�4�dǝ����	�� ���q�3������,I�0�T�2h��
���VF�4()4D�`]���� .��i�����^��
x	zͣ���t�������Vuh��v�P5�CT���`/^���t�y}�-���Ⱥ>#>5���x��⤖���_͓W��v��T�J�8h�Y�9��I_w]���Q�Hq���p����~l�Q���-��z�u�,�nݨm9�=�+|�	�hcX��ǈ\"��f�ު��:�+sr}�N��G�Q�HЙݢ䞔�yg{���z�GL%H�IB�:���d��Mi�am'�XE4*�;x���sa�Αk34�ռ�5˽;Lq��%�B����rGX��U(�^�k���SY|�D���
�\�,��3˃M�����s |��O�c<�����"U�\��+n�����|�m�[|a"���h㚿��g�P�h��;�G�.L���R>\S��s���8�Jd�$�=\�q�m��uQԔ���>�k���/�������O,4M��$.�'Y���A�`MLkJ�,�𐔎RΌ�]����9^��Wk(�"�Hy�qCt6~<�M�R��L��<PO��43500���>��k��b�	��*~M�`e�&��>y����	����蕄�D��h��PB�žC��(�����		8(\t[CF�p��E��@�	�t7���c��G�8#V�{�y�P�r�g.�ܢT#�K6��I�%2�*?�u�Km͘9Eوr����8�iT��e��1�g�@%D�&bj�p��'��FC�h�l�C�<z��:��A��T(0��KX��n�i�
�w 1n�En�d�7b��8�M��-p!�,'Sh��Q�y��
��wz`���٭�Ô���\F�W���њW����>��T��^��3w[��o��ӊ�{�e��p0,�Wy����'��-Q P 11	�k�ҥ��$?;/�Dͽ�W�ɼ�+���9�BH&W}^��Bg��˄xn�]I��.`v��Ri�5�;��mw�T�54����ڟDeZ%��#L��q,N���1���S���]����[��j[��,N��e*+�c���Ĳ\PL��FL6o@�(5�C�D�oQ�<+a�_��[�|$|���?۵���}9p	�#�A��w髸��T�\~_m�I�>�${� �>�U�g~s�,>6O� ̚"}�e�'�/&x@m� �tW�+}6<#�x=��]�d����A�L"�'��^Ig�.���=��ԉLg�<����?��Ga��6F#�+ˍhFtH�{Ya��[�I[�s����bwN*��'Z�R�ɉ:���g�y�\�1;�Z����r�AYv��ɸ�>�z26
�2�?+	��
 �a�h�WW7���Ԓ�&�6Eaa����T�I��8���q�"��2�%�=wt��GqFY�pZ ���Hi���w9C-"b��𔸚�	^Jk�EDY��l��C9,	�I�՝����\%/�����~8��ˏ��c����	]UǗ��;^E;+����bc��V;Aη��I�J���r�i�`]PY ,�̛�"�#|�'������=����S�R�ǰ��N��8z�T���.���a;��WW���,*Mu�6��$h|O
���o�����d�4��6TSq��˸imNE�7nV9�Y�U�>�	RΘ���t~���;���G�����nJ�B���b���K��o'���8����f�\>��#
�2B=�AJ�HxexՇ$գ�0Vg��9#���ˇ`V{� ���&��y�D�t�
�`�ɞ��`�0讉��>��Q�0�"��K{���(��q]%>	�(��4}NiE��cQ���e��.���ڎ`��1�l!S����ZΕ��Ө�'7!���j�ܥ��c�"�-�{G��@ GZ�lo�Nc�TŶo�cz���';�[����*)�|������XH��x/Dh\B�Eh;t�1��9Ks�~WB��&��ؐD����'�'��\qlb��D���8o#k�b�2���)@'��.sA�1���%s����b��XC�9D���S׊��P (��i�i����i��M�)N�Cc},�O�og�6�*����������,�i^��L|V�T�mt��UHeI3���Xo����r�R0�����'�W	�[�O�2����-S��$��Ʋc	I�$�tk@b�v����QKj޼���ڇH.3o6�	m�V-�tҍ�(�x9Qy0���7o(} �f�������/!�
B��4���X~;�F�w!�!�j�=��l�D�	g�=�l5��˰ ��������DXƛF���(�@/����t��о/jf`E�ǜ)�	��:�vX9�Dy +�m�Bʕز=�/tW��.k�D5��f&+�N��<�-�&:�Һ۔��3�������l4Q��SD��H�{���V(_h�	PM�d̉Cm�Ԅ���)߲�dr�e;0��U.��G����Wb�*�8s��L���xm=u�(&�ո��[��?r�6�iz}�Rb�5�{�Sh��KA��!�g5V��LPs��bm��ʽv�Բ���̇Ӭ-�j}�e���1"��ع�mΓ]�6[�|�ݲw�\}I�+��&a��c6�6��'�Dik��Q�.��0u��D�t�~�|��v�]�J�|�R+�7m��_����,,�5+���ʹ�M:q����v�b��fV[$�60ඏ�j�`5�_�a�1t!����BD���`W߃����о3�X��B�K �U1�N{*���*�,	�y2A����R���K�������M-��C�y���Bf��OTz-�O��Y��,+�z�Ż�jeH)�Ki$�O� օq�X�vө9z�F_��9�516q�^\�+��ЃK�vJ>��I�J3��t��������[�"-v�؛2��D��&m������YoU�^�W�mtD�����P_����rAƪ��sJ{�Z�= ��7lѤ�Q[F�Hp�Yz�E/з�I~AnnD;�F%�y�
"������^�{���Xۣ��s6��eý�w&b���<H?3嗹��R�/z�)��j�������SV�4q_菺Ei�O�����x��	5��4Ap��?FuZ�]+�};�9��WFdD���3YMt?���R3�7�g����Z�{/电/����yD�b���s��m7�:	���ն<������*�qVZ8�`�L^4"9���x1�j�21��O�G/
a9$Ħ~�Ĝ�;5�<�
����\����S��?����mf�<`������Oc^4˺2튶藑ѓd��V"���v~�S���+,^��h˳�)-�j1��p��� v}�5q�&rC�����Q~��|���֩p@/uH�=e	ԈYE/�C,!y�TK�F>0�]O��f=Z 5�mCK�n�|��:o�<:��x� S�V:������碩���C��C�_]m�O���G⼗5�&�4�s�q�*�W�O��pT�=u�1w�%�6��f�q26>�܎�k�`1��,�B�w�[��I���y����)A����b�:��ZkX��6���J�s�֐��� +��N35
�C
�� ��mH���F�q
��o�o�
z������px�G �Sr��L1j��f�;���'�Z�p&p� ��\q
,~�ա��Ei�P�Y�NZ��<8��~І�|.�vS�2����+l�}B�'�nfO�^��n�'}K"h #^��+|m
�Z�0r�VC�!3J�*�J��l�b9�lQZ~&�+��MJ,E�&J���{|��{w�^�]��*����~cn:�ގ�89[uW�#�ލ�ӄK?�0�Nu����LGKc� �9�#�n^�YH,�a ���?��h�����q��!�U�m ���NY;Hg�OLĐ���5���	,)q�
¼�)�����_�ӼIܕV�eȌg��������xm�l����լ'�E0NW�;;�a���v�u�8�ֱ;�cuU����<Er,�aVw�/�l����/;��=mB�-������'|���ԫ��w�/8�WW�p�5�S�s�=���)��K�����P��N�<T�&��7v���[ϡ͜N��u��R�ǌ�|��7��b�x�b��$9��M��$R⫴	�3��YY.+9u5��cS	3,`�̷1BG���j��bh�]H��TJ��2���>-�Tf�ڙ�6	f����A���\��C�x�&R��3��J�N� ����U����ҠOԄO�^���V�)�ۓ�U�K>)��&yJv��f��]�M+�ʓ�!��;�b�
��z[���CB*V���]sq��4'Ua��Ƌ�M�,�zu[�:9n�*�+�U�	03�8&m��^(�lS�N�������IN^=f��W�N>?g����I��D����=�+��V���ۨ>t���3\�����iBf��,\�3��5G�r� n06jAR���W�2W&s�.�Ӆ�����c41F�/�鴖j��ܰ<eX�D6��~��;�u�J�y�flG���.:9� �n!?�3L�`���T�DLlł5.�7ڍ*��**��>���,V�7G�M�qԕ�,�b5��b_E�.�o+�qb�����h�����T��<i����1-���#s$M}sP��nZ*m#�]��%�_aM�~��M�J�o��%����Yh��["�U<I&��N�å�oQҷ�sВ�>@toV/	7A��f���90���L�A��"�P���ɦ*Oػ�K7����oQ*�MV��Li�'��Ydõ�����jUj��?�'	xw���������[P�lz_E�dBl�X̵P�O>Z�RK�����|�3fV���2�;n@kCJ����2�����P�U	�XG?�͈��W��sAѬ�V��ԫ��E���̓�Φ���%,٥��`O56�<��P��s|]U\������0�<���~��lx,�
�g'�b�b���kd�=�S+z��[���zl�v����ׅ:>}q��i�y���nn>�6��� +@�d�v��-?����bx�!ɛ�e���ɚLN������� 6Ր�3�xs)�h
 D�@����Q7H160���w�،�`,[q��.�D�.�0���?m����/)��%�m� ;`����o����iy�z2mE�^k�o�E�-�μ�֔��{�. 8���+���'w�5G�'���?�r���=fv�WSI=}�X�wz$OP}hD?�p�	�Y�D���L���Wd�8V0T� �طs���g�$������DQ>꽃�)�k�rH�]��%��ΰ�k�\</G�T���� u�c�O;�P\�&,�Rַi�ȕ��=��g˘B�L	�Ǯ�@��%���>����3+�c�u`)%zL�N]�����ϗ�k!lu����Q�Es�Mt�i������%�o_�#��Qt�!�5ҙ����:����)�h�-����n<Py�O�g���rZ�a|_"�^�,D́������
7qba��?��4����\]I4X��Vd��9
���á�	S)�7��G�|��C`��$-��q�V* ɰ��s�Q�CL��kp[ e��"�8�][�A���8�.��P1��P�olQĄ&���@���@�r����� w!��o��(�Q�J�)l:,���p��O��	ܯ�r4-��~��|�3�$��E�c�qs���6.�R9�d�6�S���ER�4�~�	�ly'���)~�l1>Ƴ%�R�0F�d�����H�$A�Z��y�=�Ubq��A�}�8�8�O�����HA<*^�Y(��Y�ɰ�/����z{'K1��z��)PY���eV1+[��M`���W����d@V,���jR��i��m�@�"�o�	��g/�ę1<�B\���CgN�u3*�)Q��r@+�<��#�
�2��� �-`��V^+1T��;pчo���y�	7HE��	�Y�A�~��,�[��-�t��Fl����5&�i��l���ǵ ���Ԕj���s �g�s��.KҶ�=AX�B{�B�#R���:�m�5��-�'���֜w������'׽1@J�U�O�.���8Ry��Sԡ�@
|�YTuK�Pȹ�?L�9�Br*[K6� $�9��QDg� D�K�'pf����L�fQ0ǔ�S�8��6& @~%���>�D���X�5���q� ����`x�6��DH�}O��$}u-���|ֆ(�/-8�-^�-*�k����DQYY!�>�f���A1�!$Z,a� !4��!��%ҳ�!����.��-�N��:
JB��D)a����S%�8�"#��?	��.�j� ],[��8r��>0p�瑚�ݮR%��CpU���9x*K�c���Z_�yB���<�߮kZE2� X)�fד�[�0د�����Y��I���b��z�A#�*�@�C��X��N:�����|_TG����2�\�I�+a:3�cr���d���<ބ�L�3t���	��g�����[D$}X�Lq�����f��Џ��4h�'`9��A<,ɠ��G��?��8�h�(u�a|�K�U�
�`vp�S������_�����3��uj�K�S��C�w�+:+<��99��C�
O;�	�k"�����K�òq�N�U1����س,|8� �z
��M�Ɛ;!��L��1e���b1M�o�+��V��0vſ�3�1���&C����Їg;�Z�v��[�����o��3Y!�e������ ���)���a���Ƹ9KLH���Y�3��yh�9�]��â?��P]����� �.���׿�V��t���Ltpg���2��Aj^����M ��
w�C���	�CN�^k�ᆞ�9���AH�l�"�����KJ����C��6�A{�����$i�5���ͼI�`~cy������L�ɘ����-�s1ҀbgX}�s�C����&v!0rT��J.��A��;�IU~n^~��sKZ�F���5���c"+y����\���}�.'qUs6�b��&�N��au+�)Bh�(P�z*:@��<�ı3=����υ�mL�!D��S:"[��R�QTf���jG�T��zT������W�2���~U ��#��p([�^wL�>�J= ���:�(�^��B�Y�chL�+ﶤ�qI/�.����K�ݣ�-gou�fĿ��!?W�lW3s��0��$��}�x�hW$U��X}���M锍��b�{᷅�-�h�"d́|:$�J�N���+<׷t/�7?��v�0ND�N9>&�NȳXF�|Dwl�q��v�+9�1sYXLn1=s���-�d�3m������?����D�H����H�&����R�+T����j'j4�%�U�*0[�m���n���J5�� ^�n��r���b�'�	}�>��0:��@�����	pW�$��ϰ�O2-���u��z%�{��tY�v���P�U{�ۄ��{N!и��SMg�S&�[(w��j�`R-mL~��OG�qd��:B�C�xp�X}S缅|������:Ɏm�[�g�s.6z�:�Ƥ٫�b�P�F��U��Jk��+��o)�X`�������c���Nl�ݝL�ޡH1n�3>,\q��O��J�=;�iSD̓��/���0������_�m�N��}.mi��+Vh����B����!�wv�Է��� L�)"i9���$���f! ��u�������Lg�='!�8(��N�sDZ� ��>%[�gj`$Q?����Vƽ_D嚚�dd�$
AE|6�)اҠ\;s�RoŞK�^iL�c��S�.��G�Ј�莠oQ��l��K��f_Z�>u,Og9��@-Bo��xQ��s�O�Krl��;p0�7���nr�[����M�Wc�	��M������:�dM�<+�q&�0Ou�/s��*��}��k�4`m(F�!F�l�5P�%ܹ� ��c������澤�r�����(�Q	���e�>�����B�q?��޻E,0�����)�=���SZ\��^�U�)V��ٙ�ŨO�k�A��PW�b�w���mUb<��V�?�(����'.��vY �AXK_�����H�f�J7)�p~c�$�&dc���U�r0EX��nUB[��	�FQ����024�W�Qz�o�
���>���\ѐČe`�9�" ��0fK�4]�b��9��4�מ5
ߵ'{Z��R�{�o�B�)��Z����w�#���!�ܽ�N�9� ,i�v�s�Ѽ������^0y��HJd�r���� ��3f�q6������|>������Yxg�Ú��q��Cn�E�U[��"�e7.�θU�˛�G)u�ߏvw�߷���8��`�f�m+J�a�A5s����mO~�'bΤ�N��J
9~7u�&�!}@?u"̢�o�[k��p�W�H�B��]]	��Q�M��d۵3�=W_B����NZ�)ҕ��՚ʣH;�P�V�I���YW9}���r�Z�Xh!{V��d�E�'�,�Tl��8�"B�f5L��!vte���IZu�
��V*�w�
����Gf��Y!�;~.9���p�ħ9y���&+��H��d�݅��K��q%��5�Ό>�
��N+4�#���O����6#�@bR��|��T��q��`��c���0�� ��� qH�;1��M���u�XJT�dP��F�����Z�2�N{��CZ�Z7���Q8zs�������>"zœ�� �!k��J�"�Dq����9�ˀ�]u�}��e����'���2�]��1�P���=�˦���ⷦ��9D}�x��1Ѫ݄�À�c�Q�P��o�]2�΄�8��Ǻl�:���!̽S(�F{3����M=�{W<��Iq�a�<\5��)3KQ!�cl�;\��&K��Tص���Ǉv��(^ʝ7�X!Z��N;�x�$�!y�X��B�&3(�����*��,y���	�qYx=4�P-��;��1.�^��	94,`=����0�pŭ�Q��t�pg�h�<t��b��vN�_��/��x���`��;ѡ-����(�/~����9@40�� ����z�\u��
�,�)�{<�T�ic�5�d�BïaU���-����"<��%ϥO/�#L1�'GV6nQD�Ŀ�B�´�2fP|z;xL����#��������n8|`Y�cM �$	}ۿ�k�Bw����q��&����Y#N6T�3�L�:mT��0�X�d� ��^��/�A��=�;feP�u���7�K�t��^/�~0�D�_*��mYL��g��H��.!ԡ�Q����;�<�bT#[tj�*O���s)w�ˮp�ң�������Z�twH�q �P���@��b�9�9�٘�@u9
���S������a��ng;��`��O&����IW����n` ���3����`C�0v�� �����`;{���(�=q���Q�����ڛ��͚�}h�%X����,0#/�U&T��=,�*���I~X���!�8-R:��y���N�Hې���M5�*8���_4گ�L����`@툯i{�(���(i޼��.l0}���3)�^�~��~����w�� ��I��C���H&]ģ��e���D�~0�֜N�-7=�k�zOb���dp�,b����@��W5�����@�:WF:wk��v����3Ke�[��˭�J!J���hݒ��$ױ\�Q��d�4�sbW~�B��:�m�)��<�ɳ"(�^���+ICe	{2���j�����E�.E�*�<�|�c�kf�Bdf�3�m�������5�-KM�*�Jq�E�$ބ���`���g{� ��=~^3�6NDf#|?�B�-�;�pg��]����N꼰y���ջBF���/�]g�E��{P�)Gy��.�,�`�W�c�ݤ\�glf;{"񓏺˳�r��b�ò�7v�$#���0̨��-�&���g7p hU��/)���+)l�+ZW.a �JI ��s�d[7�<�z!4X��O	�Q	���[�����^�V͙�x� �*a�� Ү�uJ�g�*1��	**�� ��!��7�*Z�Gt���C�O��Pτ΂m���ui6�a�����Tt�Pj-�ဈwW�rJ���fN�l�A�ȣmIM���A�"t&�A`37C�Q((�?Q zJ҄��]���QJ�Fi�vXMq�g�����(�ⵌ&1�6qG�>#�͟���Ĩ�H�k���r,�g7��?i��hv>�H�37�	L�@�%�v��n�adz}�Y����,c��ynE��X�@_J�p�&�i�,0�&��Ii��?`�~�qk�e�h�K�v��I�[_r��Ea���N�E���]��'��"5�q��Иz�]�l7E�sf��'��Kk�Bj�Fcz���c�a[��E.{�/0�����*�9j��А	�J�>�"��xMj����iK%	j�S�%QW��]I�1�d�S����oՅ�JI����A_�o�F'����d�Ŏ����!�*�����%F�9�XT�<��oJ�8��%���3ɗ��ᒅ����%o�x��
ᷙC��穠�����d��G�e���7R�����p�G8��,����o�'{�b{p��i��fQEB�Q��[��nc{']��J�bՀE E�Pc0o�T���*�P� "�c�.���'�-*)0�(,	��߹�?)>�k���:�. ���x�W/���(F��6ȍ̟1P�V~ 7�k��m5Y�K���7e�����pWF��	��K�>[��	�)��N���DL�)S~���'c�Yū��~�xz�9Ϩd�^�B�ƻ$�(�\ͺ~���~<��A_���B�ҡ��OrP��`6 �v&:c�Il�j���oZ������}�����y��=LfJ�X�}{�e�6��͑[�Cc�O�Z
��s���٘��bV�0y�(��r� =m���
���Gh?S�`�*�c{�r��t�4��4�gJ�n�m��d8�Pc	���L]<�޺��������X���n����V⡍V�"�w������@��<t�W��1u�����J�#����?P����$�п�m[�4e���	����"�ٚ�o���R`���>�֣d��'+��u�Oi2�7�lv�V۳E��\��[�(����DS6�(V�Կq�F+����#�1����.�/��Ό[1O��~=��X�|���d��I����b��Y��u�1R�"��i��Ʋ7I�;�C|!M�6���8�q��L�ҋ�|0jO]��P���~�b�B)���/t�$rz�!Xd�Ώ����p�
r��x���lG� I_�n�p���_�S[1
����v������Lf�����3_F���T�i����u���*�Mޟ�{eL�0����Vj\�c�.�pp5��~�Bsw��6ty�X�KR4W@�d��q�k�
Bn ��v^�\ZX{���]���V�� �T֗�Sy�?pƪ��l���U��We|7�;��OҲ���zB&$�yS ��F�6���j]��=�$(ᔜ�m����gn�z3?������j*6�6f���Lݡ�+,~�&f��A���	A�<�J_�L���M���w*cwtg��ށ�ĺ�,栩TEF�1�Վ���l�\�&��̎p^h�&�&)zy���}-HҾ��n)a(�^t����xx��\�/c�i��ͩ]��BZ��ͩ��(����*�H�����Vў� �x9z-��^(�{����(��[�v�#R.A�}x$=�[�V�Z�r?���bY�.�.����f(��K�]?y//�ƕ'�B�{�Z$;?X��4����)�1��V��9Jw`��N�,^�J�6���k��,x�;���p|�\k%$�x��\z����H�N��?|#�@�	�lo�>�����5+/�HU^vå)m'�V&�`[I*TM֐\[$����8@*3`���ll3zr�*��}(�w"�O�4�;�2O/�r�Ĩh�T��(�u�=,[�>����mYI�ޅ�<O�0[b��a^6�߁��%��'�Z���O{�R�L��E���LMl	�)�(�����||)!��H������H%�J���u�y�M�L�4��ؽ4.��G��1ns�N��)Ͽ�5�L� N� ��7�]��#���7��F2P�L��"�PiG�>ʒq҅��T����Λ�B~���ϛ���U����(7Q�¦�R���_Fe�ԛ�.jWҜ/��m�<ҫ�o�Wz�;0�/x,�"�fS@��e�	��m�������~S�v����, �24�S���4,�J�>u�'o�M���i"��p
�N�gOK�/�̈u���`���ė�5{�!1��껼���Uz�ߎ�s'ο�dp�Jxi�L+�6�R<��>������~id�ڐbv�[��b�N˫Ah���?gp)0QB�a_lR���en��uZ�C�tzq���o%
�.�-�qE�wÊ�K�F�T:HK��)Y+�Rm�mĮ����#�8�H
�؇�k%��|ʡ�Y-��ܚH���h��rbTfܗ�
)ʇz&G�"��BB�n��!��1�Ŋ>�������P���^#WP���E,~�]u��𛘪�e��%`O	~G�h��[�F0������Uf��u
��9��r����8��7�S�g}y����ʆj�kX�<�C��]�g
i>C2�C�搬nf��?�a�?���U�����>��jk����Ff��H[X���,������H�N{@���rIe��S��NsA!���φO%S4�Z��ǹ�#f���S�%Y�`�ak����a�ηG����\��q�lٌ(M��Ae��������ᘚ�s�ܢ8���7B���5af����h�8�C�VߏX��N�z�V�1����������[��~5����>�)�˳i0��J�y���b�?��z��z�GpZ���8��/f|�f�'Tt��6LB3�!����y������"�q�"ȱƊC�U;��)YMR�@�*π1-B���ݜ�A!V[=�/R�b0���u��H�NB�F�bؒo6	�ěU�����l~��:��.�h�Y(ј�0��f>��[K��r�A�O�ٱ�m�w<�T�-(���I�_�O���a��[��Q����z����o��^��(]�M���BHZ'�IE0��{��o�X�e;S�x���nŗ��"'����M�4 �mx�?�F�|�����D���m)�e�f��:����m@�ۚH����r:=]��G��W�0;��~���b����Jo��-Ƙp�`/�}��d^�ٸ�A��6�WԕLh��"8o
���m?�]@��_dE2;��[���Cn�A�
i^UH�t��!��ţR�%Z�G��rQ$;xQ����L���t�GБ���ۧ/��iY���koPp!�X�)C4�X�)j�����Kx���oK}nZ~ȋq��L�A�$�C�*mX�Ԣ
m^/x��'��MM��4��};6U��zDg️'��23�os��_�� �A�P���b�\�*⌵[cv;�~��?q=�
�����>`��K��n��#c�"��~~�����,+�y�{�Ϻ^��R�xdm���@?G��YF����JO�����gAIňck��k 1Cl�����+%{4��;�bByznwyyS��f�m{���>�h�:ۛM�,ޱ�ws�������t"�:�6�=���n���`���P䉘/���,73dC3�����y!�vex���W6�u Q%�(	�b��H
�[��MӜ<�P�R%N�(**���<�R�A���o���2������ӄ�_��(�*��H0pUY������ɜ	K�ê�cK���"L?� ��!B��h�@�A9��3��p�}=�(,Jȕ#p��F�W�n������_�W��ivE+N��%��,���OnB�]���g��R���;���0��اJI�FĉB
$l��A/�i)8��ϟ��Q�`�fB�*�id.��N����'��O�5�]B��cD1��>�o��nͫY|͐�o��T���=�>=���nK�?(��o�8�c���܆6�ӫ��
����Ld�u���f#2㼔���|1�4�K�i�z���B����_m+�����la��t�O-���*��\6���o�g۪�f�ʍ�'�}%a�"�K�8Ʈbk��z_6�)��4J����ċ��.��^�ʚ<��O1�n���K��� ��9���i�s|nz��8ұ��9�:�̱"���-�Պ��,����ӄ6_3_�KI�ga��0��h�hw��>�n����t���T'7�n��Y��U.?�����F���yeb�x���e}��j(x��_s%m����h���KM_N!�؛_�8,H��������s�+�LD���]�4%��4�#Ur�y��;ّ��o����؃��2٧�+腨�&ܕ<���>�VI79q�E`����Y	�(�I��ʫ~%�e�1�:�cݘ͏��*�Cb�Ũ0�_��g�_����* �T�>��&�͹\P�l(�#)L]H��2��sM���س�t�O���Hy���#d���n���f�x��+����D^��(q�|MP��s��ҙ�����}�3z(��7��:P�4mA?7�g��H��"sr�)"�¸2������0��3��qV��ռ%�v��O��(=!o�)c!�=����_�;��8�	��V�Q�1��*~�~+��k�s�ͻ,�z�t��[hQ��xe�6f���M�K[m��J����n~T_F�-�h����h�=��[yX�6�f�^�XZЀ������B�J��\�|-��	V2��}�zP���Q�	�4��^�[U��\4oǆ ��M�'�,?.J���
V �- R%e�B��R1Zʖ=���&\�GZ��,�����{�����z���1G8w�y|�H�"9��;�5"�B]QY8?/�(���"�?�:fB��9.Q�u<9ڧ�&'����d�I���|��\9 P�=���b���t%F0�@��?{s�ہ��KQ��;aDy6�^rcC��?�ǁh5FA�2y�:�lLH���(���6/�>�	�?U����|�C8T+�����9�acU�p��l��F���e��8�n��,V�ٓ�;Q@@�
�P)�H#;�ݱM���R�W�
����a�I��)U̳��	dc��J��9��,�[�c��z"d��mһ�DM(��'h���ixM�pK�.�
<�K��D�xE5@�jN��GZ����g���r������=r4��+~����@�lw�U Rm0O=D�<�ы������Nx��L�xk鼀|�lvo��X�.��萺�El�s!폢۟�e�A+@��� 8�a��ٝ�ύ8pq�|7���̕������F��ceE�5F;;$��"����Q_��ԏ��|�7�8e@eg<M��e�'�*6��v�i���=�
h�g��[��Bj�-��k�;2��ؤ�
tqd2���9aH�$�N�B�ɝ4b{J$������TA��u��RUzT�D4���'�s���M�hvr�Z�"�:�R��.V��A��$�)̘��j����"-2c���߹<B,[g�;��z֌��Q@�lv6x�"r]�3�kM�?��a��ҁ#��V'n�C��6�#�ɂ͓�]�EfŸ�r���>�f7�p��}�U��/��k.�����öh������m%����!}�qZn�@05���t@o���v4��-lD���d�WĆѮ�T����*�Z� ?�S�t�?�����./J������UN���Wn	0���G���;5����\x��Dj��{u��³�6�P�|��>.���X�b` .�|x���
�Wm�'�߁kR��#��1�ER�¶x�;��bﰔ�C��p�l�Me�sb�x��_wr��z�iv=L�ԭnX�4\$�DK�^k=�M�VSH||��\��k�̵K��0c��%��v��������}�5�ퟡ���v����tě�
p�R|f��4�7��p��E*B�1�X�cy�,q���90��D`[�J�ݒ�W�$3�u�!�N����m����,g�y�ă�p쮴�w�����j�Ŧ���m�?��$��B�u�Rh���y0$���.��;�e)܄�ڥ엦��U��a��Ȱ�1
[iL�ǻ�P^6L-����:��J� �t#�:u{YW��c�[��׵�ůs����r��H�;��s'����Nk�!w��jYM���{W7VJ�8��d0��~+cf%�^NY�5��dE��Y~�,b*�ڴ�K���`�l�+v�}�s����ҋ�$�UQ=�uT�*B��\����,�_n�P��^�"����D�G��8u�#��5�"I�-��V���I���-���^���ewTKHNw�R�|ȭu*O�z�7k���5~9��p�.Nއua瑽[��*7�gw_�3�<��3�X��FKt�q�o�d*���tp��{�ɯ��x`������q�B�tW�W���*AI�jc�[�mQ�k*�p���/����Ss	i����_ip����aF����֝ �j��d��hτn�^�)z�Wğe�C���nH�S��C�W�O��x���n.yNC��zE,(����D��V{���Ň��J%	ݗ���:��+r����m.��my�(�jU͌������c�J�͔�n �XbU�a�ϙ�y@س���M���M��O*'�������6�i�\&��3i�<R�FHf�X�~
b�%�M�0,\�������ˮ�ݍ����S3�
�" hI�Ɗy�aˋN�
"ͺ� `�g�ϟ `�
� ������F�mJ,�+�a����;e�3��@C@��1E1M�*b�+I>��j���|H�k3u��P�)���T&X�����H^]q#D���(����OY�x�QG��{)�
�?��!�= ��A�3ha���ɣ1��O���ްf�[&znfKF��m_������wwB�U�o�N�輿(Tn�i��+t��R�hN[�λ�%�5$���U�-�+_	��V����S���������9�X_�Vch��J��Ґ2��v"�M#^H�	e�	��=Z��� ���'9\i��b��5R��x����k�,8�+�"ws⋍�Ç�25��zݘp�v�"�DՌp�wQ��G�>H�!��a���Ɂ^��k���P��؉��J�!�'�Nc;�OS�v%Q�;�(�0sk�����[0 ���Y3[5��r�.(�^U�J¢. �>}v�]89�ߗ�?�����T��{A�1���^�;�猥�.���k�E��2j\��2�:��=�ҧ�gPH ��|���{��]���bA+OW�T�� ����lj�S��� y���BY�]i��n)���5m��:�U�35��^W?��5n�����bp��fh.<���A�U��Q���^�@ƣ���U�k�*!���} �d���<�v�D�v�AD���}d@������6���o@�'�"�t���5���[��aVHݘ��b1�A��X�Kh�2�d��$���=�u�ki��*��cMZ�c���F�p��ifK-��B"w?XB��|_2_!�t�`��$@�
��M�3���@$��8���uh۫�R�ޖ�^A;E��UK��Ka
�ֆ}�kƄpf��ߘڴ1D��"[1͌�ᬊA(�Z��$��
�R�����ƷVһ�O<Ɇ���p �6i�l�˭D���lք^�������OgK�B�C��@��O�}�1Y�-�יP��?�-A+��0��b�I�=	�!��\�>��/À��3EzA���겾�����c�|�Ko3�g�	VD���_d#�%��՞��=��|�LbS��[F��ٞ�s�'�8�����cٞ�o��M(o��h�+���C=f},mLΤ�v�#lX-g=_���ʴ�nO�H�͑Ȇ���!f~V�"G��v=DC�[8gS��Q�Le��u�$�Y��h'�K�p����8w���6���\��h�GF?�u�L�7W�P�����gI��~���yt��������a�*���v{��?Z�0�r��x!o�b�}��E8���\"�"�BQ���dɔ��?���%]J[3�q`�\��D�.~,������ ����W����?N� 5��t��4�l�3"
�dIC**�>����H����'<�4\�A=�!B�u�'	]�3Q����x�>�����-l#K�)H�,��T�E�6q���?$�`���h�2�����ؽ�����u�4I^/6�3�������J�v���X��\"gj}�M�Y���bx@���$�[p����l��N���`$�-m��4N�8aS��k~�~ :L�ih&�8�#\����WJW�)�&�3dee�Y1W�E�~�4��Av��OMxN�[�ehF�&۹���7�P��O:O{��V�J����~�v�����,[�`�S�"y��T��!z�߽m�q��qA�8O��I����ʻL����m@H�>1�ŗ7��{R_8�5x�a��z��uW1Zb�U��B=��i�fо/���0��X'��d��WcS�=CS��}9K<~�޽��XJ��E�K _�l���j���W��pCS}��k-y#-&}:8�0+�7��s�4��>C	_�*r<'"]z>)>ʛ��:(���8�eV�G��aWaXHv�z�_<�H��3�q����7a@fp���EX&��l�f�G��fx�S�m5�fʚ��lt����0�2�����l֔����![�~��l��Aa;ԩ��Jsn��y�%���~g�5�ǒ	����7�<���[ֿ�"r��o$�~�h_r4�P0�7��_����w������u����*:��x�#Ǩ~�wAr3�g���!e}fj��m(M1� Zĉ�L�(�@>�`�D�5��7��r�0E1��z7�\�m�|��{a �d�J���l� �5��oB�K<�x����VP���H�f��pH0�<�ٺ�b)��縿�0��d��k���S�«���ӿ�Y����B�=�$��6[��c
z��8S����wB8��	׼���H��v*�M�I�V����J+�SW�Q^��&�F���Վ���-Y�� h����_o(.v��� q�g.�a���k�R[.GN,��&�t�[D�g3~&Y����fvj�8����b7�
��F�um�FJ��2b��a��^Q6V�Y��Af��)#;�)T�����&=�>X�����fyA��~�>�$��꣼�q1�Úd�v�9�~K\��F�TN'o5��[��� ��^��f �ʇ���o�TWA�j�1"���� -K;5�$��F��i)�CI�jB��'eY���ׅ(,�U�;n�8?l�y��1=@r9�� �lm�)[6�c�8�@&�NNqؒޥ�VI�E�ͤ���FlLl�9%�>
1s2A�A���MJ�"�wZ)>�AD�4Y��8����w�\6��B���]� q3 �~��`�.�{qgx��2���(�Gu#��4�Ջ{3����ї����ǘ�M�^2���ma���ac��}��{�$O�[���QZ[^=R~�C�l�jy�i����~��I���5�����r'�a`�B�\������=��.��G,�&�T1/~K6	�j�v�V�5��sK�&ޕ���-�<P�P
��� ��]	���E�>6�&���t�e0�v���Ŧyt�UPP7�?=ɛ6��Z���FB�]P����D�ua�ѓ���Q�>1Ƌ�a&�w �(�;�S��WF6癏����?-{�0{ʚ��X�Z��36w�tb�Ip�Q� *��!�����4'K�-�ѕ�6�b��'Z($ϝ�<��g���(��r��D5�&0<�?����s���"�(��߃Y���φ$F�5Y
<��gK��^[Z�q%�p	b�&�@�Cм	���^u2�`�-{ <$y���6>�o?��v���tlWS:���v�v-х�փ{Ox&�T��vBH$vLӲ��KJ����ciש�}��SB��ų]�H]�7~>o�l?+GE�>y_���t"�!��r���tszY��߫M���e#�kx��Yk{��J9�,�US�6��}92#�Z�2���x�lmx6%��@>���u5(��;�ݏC(rق���(��i��شV��}���c~�GS>�t��%���>K=����{�k��|(  ����f*�V��F��(#��Iri�^!Io$Jv�;S���nDf��e#,E�f����|j�Εm�o,�k�嫭�H8��%��h�ˬ$��]eJF^�Fi�b�2=���U�c��~���G�	�认H���,M��z���Lm���QG�ۓ�8�=�Ի��	b����-�ȫ��.}�3�d�LO��} 2:ɣL:��4�;��v,8�Y���[y-���*���ғe�L ��.�rͶ�ߵ��D�g�c��Hb�r�	��ܼx�ī��~0X:vF����g�۵�qR�.�mH�_=z������Tό>i|�Rq���c�v����l`���{�?�F��.ıx�ȵV�թ�=u`)�����k_(��������2'�$�/��rC2֎Dn&�>rN1F���Wg��zz�k��顜%�����5����&Ž���p|z�:#ʚ�-�B���h����HKA|zl)�- Kn����;D�]��^"iiH���D4���ʜ�{��9�➸ć�{���51������XW�r ���{Fl�xřs��S��?&S򣟭�99.�L,isǊ�R�/p�q:};�P�HK�Xk���J,I���lds����R�c�Q6m:&i��HI����܃%��f��F@S���7��DYP�7~E�o��K/���w'h��^	�p�X�S��'"�?c��V���*j�����c#_�
��v�`� ��ط�WbG��k�P����?r�h�@ot�_2cϯ3Ϭ̭����ӣ�H ,��^��'dkU�2u�RLWx�g�3t�Čƣ�z���6�ns��pQf���"Ҧ���k��H�'�M�-_�{���%"�j��[�6���!��/R�����x.�a���E�:U���iPA����L@*�w�h����������
���L�w����haο��eH1ޢS����|���x�ڬ'��2KQ<�A~O�@X3��d%�f#�?��4�*jbP ��3��Q���Y�� �m> ]B�6c�iĦv��~��diᠴ	/��R����	�I#6����(-�9�?�=M�r'yv�5[�3��'}�)�$���#p1m@XV?�T��.�����Ilt���� �
;�Y������e}��⌗Ą���GC��`Fo��Z�٦�ǑEE�&c�&���o�?�u�<�0z�%�I�,t;��7�^K��u}�=J�ԏ����M"ٶV�#+���`� 婭b.��t�)v E�nz�K���t�z.���A/as�]���6~���)ZO8T��F}�Z	d;��uq����ә`���r����U�$���� W�Z�Y�g�;�,j�;f�q�ˤ�
gx�N3o�3�:rn2n�m������ĩkB���8�^�ꮷ<������;a;",SdlE6��ձ=P���b�z���
,�(y��B�Ou���o��((���T���9���G�	���]i�ϭӏ��X�I!)��co�-�v}�-�1��BĦ�6;)�"��y��1@����ےk^�ri�ׁ���������Z}uG���6DC�zƼ��ԶD�����ϝ��/�����V1�mb]���o���3d�:Tg�|V�Q!��y��4fg�܎<�\���\�?^}��,|���<m3F�7in�0���U�,!�	��Y����0�qبB�d����5�9i#o�:��IL�;�Uh%�Ǖ˩|��_���7��/��0GK�B�����o��0D�>t���z��9�!p١,�>'�f储�]�ᖦ������4�k�F�3�jH�B��k� ���6��?/S����4{]}����^�q�6"