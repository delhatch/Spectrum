-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K4o9lRMXzU4IGDin3QPjQHPPXNqBvZxrs4M8L9j9X8Jzeec69/btGIjY/WoST0O0S5MEr5nNpLh2
/NKECej42m1iQqrHCCWmSSNSfMrECvWWHz3xGXkKBB+MH8jP7/58goL6eEFyvTzCjmN84EoSLiTP
2uPgELru6NgLLOrV9KTVb5SdhhpywPHcPmpoDpwF/P0TA24CZOTZ1HO/nZuwF28Tfj3UQ1vVY35F
FvfsufOJMBY1BoF1TI5lew/Fdb/A/R+vyfuE0NR3TIJzdEbguXukaXW0mZ7orWPWPBeRjPCNqWj3
ijqlNCBuMhCWA2aeoi14UO6EnZcNI5wJpQUyjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
uSPVNcpFt7pmTCVSHmAATyGyNb6RTy6WDa5fFFdV3W3YS0VwTuIlz9Nb4kriAkdT051LeZS9ERN/
0CDnS3FY64iHsuanCWnq4b/HgLInnEl1u8oJFAxv8Q2rodsoenLIR8njSA2LovXLTvKNztAWQ/RJ
BMEb1zHnPD2S9ep83rvNye+vLP/iDc2rHmVrRMqs8pfZNv1VzH2aH54dXK82W1mGhz8OGccvGHxx
5Ove6pbHzXErKyBg2HQSa8A/ihUF2R0xYftCESceKrhhISwkYvzpIy4/zgPMiytqps66zSSr+Psw
OIpBz2SGp16NsPxQs/gzufC9CapeuMur+n9FAPTeI0upJ4iXNTBzezGYKVNo2DC9lDHx/2xNZ72K
ROvLbSG5KMfUz+fAWl3Hn8UTfJpgCVva7NLkusqhpKaIGzni6800oWvZNK4xw9rzENL9XglUhp1R
HpC8TU/YB0c2xDOlFyI5UNaLbCe5DJjVEsGvUpQpndwhGxwQoG6G4x3kY14jbSKbQtno5kKxiYXj
SuMc3B1n9GqvFsGppqhWFu7c/tV31/iK8r853iyZ43khPinkyXPcXxI2OX48Q8iZFo5nt+LYbYre
vSCkvxVUf9d++inKNhxUBHXFUxDcUm4jKrRbJk3/ZpSBEh3NA3OZVWRKkus/hHDZfOwWeOWYX3B+
hqrBqjSInUJspzZUl1YNCg25wScYvFQOHCPVEFN+80Dj0lMkor9AwltJAyv62cjqYLwmq9RP0+rR
6wSoU4muAhWu1DC55NtvnCASCI98iJ3x5scDSx52NuoXIae59Ana/WHz+hHQe7FMUvZAGFgAqyN1
0C5ZHhvIkg8mhjAosCPORnj93jXjhMpui38/o0HraUwhgsL8UmuBYWczgfwBP/6HQXP51Xxizta/
oibEh92SOW1PU0uvvmoCMIP5+y1YPVOavhQ5qNHAsjtXi1ZtA3QSl9ZXc7HaQPbgaWjXZVHCa7bT
zWCrJs0LxWWniMKn47O6kikyoMxE2KkEU2XY68XgIBDc9DBtzUFMJQgSfQwuYlUd1romSH5K4VWg
ASytzIkVisLesnh+mlWUK0wnk6Eb/Zq+dO5q3F3HJ4j2IhTeb2BmRZhMjpIf2+h0cRmq4eEdElii
l0jBbvL1bhOvxp7FMV6CIS509XpF+EhY5NYl1Gljn1AFn5HN4b3ENeKonBgJxXtzrh3f6TDLMx91
jz0rDp5XqD+b3IzqDpXZzjOLDaI+pp8U2sYZ7zj6IbPgMmKTVz6dDrbb7npGOjqC7wIGtRvUni0i
TfpBZUniGxUhKjyd+nySq0NOSHT89/VUHoRW3KsfYvQ+rusWb6BiJnr2136XnD8X3TQQEIMRAL8y
cPJFWmuhs3d8skaHCFCarHdI+R4tACdDxK6BYP07XAcRXmNueN000WmkOP3U4vRKZI/GRfM7XBi/
MOsZohQzGePE+lDRCEfT0gDOQgjFr+/R7f8fuGQ4k+okj+rNrWmttPjKPgd/5jquDiqhj6rLLxyF
0tma8hssCq8Wc07ARMc75HUPy9PqV6QbfMrb3HLx1MKPJtEtIlJ+K5bcYsseT3umxoyM+NixNaFz
DGm/Rr/Mwt6nCJYiGoJc13yi1OiWuXOFGM6eeYa/YeVwx61+X+759X32HF/DZ8pKKn7QoyTXKY7k
tcP8X1owALdtXU6vj00DKtVtklsfurnpIStaZKAQK6VYn+7IY0K32aiSnCWlKixSayOpk6YWxT81
bbXA5M0lNO+Y9aNG7Z8vCcyfwy3SrlcQW7roMrc9/sma7h8PaCHv7N0EwRyuLxBAaHAdVluLiExx
RvlZcIwfOpPyAPHBYiuVcQmRvBjOj/F3KYTJ0uZGWM+LMO7KS7tZu6Lrp8nEisTxz+qP8/ugepbZ
lomubAqkYuvyktXJXNwDvT3D7oCcA7xoSqw/UPUSQMKiU1P/myFgpdS4g/TDNK9RGjvZscqsi6C4
DYDsYhWks+pB5XDLBJf08HMiwtvvoVV33HcpX5Xm1cu1n5GHoCNWzpB7ykAi4Dp0u2JysdVJbI4/
r9DpUZzcuKyzTDNZGVKeL8PKu+5n4N+6osPWYynC0kJc//3kaZ4fey0g3VvkqsC11GtedsR5Vc8h
0s89udYVee6cJiNlSDaeXZqbeIO4icioUVEPrHz3boUUiapOtMiu0S7+iuB0ClVfhSz0zunAnBKa
ZKfuJjclk5QEvrWI2ETvsuJPynHIrBlD7eSHLI62tQ3dK1boh1wTpIDljx0++9uhSqfISmmwIb/V
9PYQvX8+86RcRH6LICbf2ivOERIetoYtqsPqN/eHDYj042bqwZHGfdwE9hGJ/wQ7tAj3JkSgX8go
uqTx+dDsP4OYNGa5IZI7QqwqO0Y/iLiVZWCY6pNUSTT8OhRdA6dGqJ9r5ib9q9rhZM4ZDSb9Ds8F
d0ZdjJYmNEnPU6Sf6PFLZo0Ti0z+8qVPIsWjMAQSQNFLNpjUrXjBqXQ6EfLVjovbOlnwMnXcb0AP
0noBlZxOxvK+GynDJGk+vqXfWt5xJn7rr0byTjdkO1AGJT2I+SEGwpVO5wiIDUc9a5AG/yrtb/LG
X2yeSiYM0Jkui1Q9Eao/JKagvx2xhg7tlgmYL7OmAxY5+v9J3QcrWT/Z1nigm9MBLuAYBrg9npAP
Vmckwt7yBRk061df/c1YxSaDCF1mQGnkd3y8GHgusitM8yFOXwmEmRLJWwyFetEefBsLTH2CELSW
VPHPWc+0py14Xu4nlrY4PY47Xd43YvS4sUq3ydfuwNbBmoLHjd6z68ddfQOV5w6ylnP+Vqb9xiaY
6pazOJ77EThGnzHKFR5o4HxD8PJlutVdH4gLka7c738KJVAQr72UTa8j243c/tEKOme5+9yovbKN
KKGxbOgV8Tiy63z83vaLKY0E+oVTMhV3i6EPNoD9B9hJgJpYihDgjBqGYbIW+UzqEIByrRIqHbr2
6QhA2tz4LS+2bsaNmmIUBwfaBDJM+HOBEcoNM2U7JEP538cTOlEsxwFqyttAliMzGxoZcaeZfGTD
z/D50Lxuxzq6tlYJyjqVeYygAJEFOBtf/XnLRWub1/us3zPzxA8VQyhyKTcVOUHnbgXScfzJJM5T
QtbJnkT7O0JtkgN7p+CJZxZq0tJjYK6mFO6ItlmFF/m4nNSqsNF35/3m1EJVcFgFHpGFrr1MJSC5
l+mHgooanNpmCdh9opkcDaHddqge8odR7mN4m0SPHdPYhf81aa26GrpP2pew2Z1i6rHaF8N4tKb0
brmrBDGPI7auqoqa/Gg2AwcUbjga64x0AlK6WPNvYV37pujzenp2wFghxBmjUjD+0rPyTaxiYdU0
7Qa4VZt3htqujKljWKdzSzBzIAcwI/2c+100+/qY6Fqemu6uIxbcZXAQgIxsMxsT3q9FUouLGwgq
Y47nhFXwoD5Q+0bljEvOPhTcYTrt60gXhl3a7Fo48B8Yyit2nLNIkItMswDLC7Vsa7ICNpuuwtiI
KRI+/k6zxOM/mBdCP85sud3jPctPeiiNhUPcpSb7ol0h/qw3curuOJgagL+IbWrUuH4K+twBWtXp
K6+DrnAtSedieQZfL3Up5KonSRjhnVZRFrcR503OOXgvFobF6MyKbDdZvcaDCsfzdfk+tjOzAP7X
eFjgoe7nHyitBM9ZySfTMLLPZ9GHv1hnUgLUb9Qy1wzzdj1TV46LCYIvFILLT1GKVR6ZNg0VcYrr
NKBD7voveyUNFW9g3YiVjxSWM/8Ad/st/9kDjry8Ts+W0ZO26qVNBfspk47caqWFjFA8MJ5Hdkjy
SXX2fpPFPaB5gITk9D6d5YFLorA8ehHiTOq4h3DADFDSknrpZySI9kr+uwIv7UtYDdm7YGa3ALfv
0ES/bSBDgW9hELV98K+RsblmFX5wp/SpIlTHLyH3zRzs63iB7aBV3qKEeIzsoRQrdBa07G2rC116
3+0Pf5ft2IFw8DMNgydkvR0nkto7NJ5KVI5eq//OX1d1zxKQVRtl2Yn8QGrMTdYPCMbZASGhCvfZ
KCFS/SFH8CWBdN1X5vGnRGu80ZdDiXmehxeqKI3bCIqDFDSl4ZtnhV2Qc0J2p50o6+3RA6NRSUcv
1xbQTsj3Yr/ZVRFbCl9RWyEw1mzVJ7FVKaZ/qF9IJsPGLDlfl6dDNzZS8hkbPqSjr8DXLG0K7N11
QXZN067X4l9fqL0hp/RQNv9JO6fpo0JkNiNr5gObXU5E6Qw+JP/CZjLeFJ5aCa2dbtpcKsgb27Of
/F6eN6XwLmh8oldoG8WbNVDFQYY1jewMxK83QN0vRJeUOh6NjimU5Ur8Xb+fi2ReE0z1PuoBaxHI
O8Eb5dCOLv5ul8w3m9aAZ7FPuObRnSUrVs8IfKIvaZOnxFcwM+XtBel6Q0l0El+/0wkWGJp3n1tU
+/dV2h8ZGiuzzv4aaA127JMfNCHUErMUAwGcG6uG7FpCpHO9Wdg5Q/v/xmb5ltgHo9T4IK7Gj1rb
lWddgulyWXJTlLIP2BqCJ358BXTTePUkUhJeHuGvPPTS+lNbc3PExpEf0RwkEh12YRiUnfPuoaca
Q/vE8LjRp9jocpniQulTP5yPUkC/jMLLEwoI4BlETnSkbfU3UXBBnFkhTVEwMgWcmAd87xzXI4WC
ExuPNOJS1etYWv/QdSoNlerXm1hX7Q40eK0ybIXlSwA9pl6gsjLom19mNCkn0rdTI1qGUCStfDGt
0llxysqRoerjuo19mVHumJQCH0Ofnmkmchtue7FHSl4IV9sWfztaTEwDPQ0x0ljp1R5dytw0UfbD
5uqcXyRm4pbQ2NSKK+xtM0WFCvbvjPDIMfpLPZq6abH3eR7bcmFdNxHEzxE1JF+6Ig+u98jmJLeW
WVKGPgGiezBNcH+b1rVWeSd7484WaCDGxD32Ra/f2jsv8Gvcm/8OGtWj+IIK36tA82A5ODDXECRN
FvzZkyV0ACQtHyypp6Un54NzcX/R5gS2MzvEtHrVmoCVRtpfd3kEXl2ynoKFYvf7cQOnZpwadFyb
Po3RItWQEPXHGr4z89soXy2DMYjmk5fH1igTrSW2K6w4DDjWEw7RnYeq+myKCYj6ddq6GNKwRpN1
R8NS+R29IDFwMxu5UPFvPlb40YdE8Ye1aqObMVsEBWbiLH2QwycAu0BWC2L5FBiNsJlsqkIgH8J+
LtyMP+599k+TDqGb1W5pNTzboXF1XbfUwIqzy6W9ZGs03Q6jsFH2MGa8NEokuqR1s2eQI6SDGqht
6A6w2sTDLHVW4th/6ktLxRE6BPLI8e8Bx8JaMHflK9sX9E5ylZcZmy/VZLcMyNDGFxmbQxy7E0k7
P9xaFL+ZaCEVqVEx1DcUGMXGpEfUPo2IfAfpamoqU3C05IiRKyNRJ37cH8mibRpDhP0XXi4t3Px7
04Md4SGKEcCeCE2bYiojKTvUEgg8hEEYRlbKy011mSRNKFnhuVFwVdwq6NdjgHB9tUrT3mGCusfM
+Dcpt6YALg5NzQaPlKt+rP+Bxyk7APeRt+Uw8R/UYfaYkMg6UCpwTisvRXLKYMpvcnyTwlzIUtkF
PbRgk3DLhMbLHZAS/+X0ziSpocugZvYbLuin52Pcx+2i1wwfzXCVTv+LJWESAIwwwIqolU9D+PJX
CoymXptACQMDOEtbW/i+oRxjOzuN/vxigVqNw5fEcR5r8LcmcaS//EJpMXr2MbYkdztiZuxNVQaF
nhBCocR5RBlobSGjV5cxylsmiRxqceaFyCoRS605KKm76t8qVjELhL4mpBFTkMB4X+URwZxtvdKr
Y9fYTxOOWYAgO6JY7m7pcNS5sMc5H6rAXVuL8iCiQ4DzZ6JYXs5fK4VkKSCIcWr4+JcKOYuIwArP
9myPIpTyP3Vi+k5SqhX38L4pr0Vrcyg7IcfJf2TWyGJW4ub5O8qBSrrkkkwR4AZXqwhbCkR4dAp8
xn5Y01EXdVgyo/gsUrh11UgYEgGsFjYR2KBJ6gP9P5AV/wJSnm6G1Oz/VCLXI3VGDgXXAABu6qdh
wisf1W+ZJ2tnN3dETY8jefRsDKy4SWviNDg1MTfz3SdRACdC6M5tz8SWqUreRI15eoRCWMoKn45s
QkulafSa8ajiDUqlBsCZx2UDcRpqaVyxfVsoWJGxPLkAvkWsUPdFkcytB4CgSMagzydf9bb76Few
4wjcf8CxLtVkFA5ETsUxKWWkIb4yHJOrl3fApE4PMuMiQsBG+quYyMPDyARlVpYMx+kRUCKWbnsN
CV1OR/I438fm/PgfEZGyjN8QVr+jhA1ioqaeX6HIyMWARTqwOdK7rJNm2y6hdZwqm/yeq9tltW+Z
6pxAdIqnELNwMOYPPdwUUwbDsAYGOMdf0wQ0s0t0wsmf/xjrzHWeEAy3+KcZVQ+ah7OHjMCarMXC
vxNWhoe9+jo4/yxB5u/gyd7aTuLAHBCqvr/yPiVlxid+4/oWrsOyg+cDeR5B03zGJ7UmGn6seE6c
0kvp2dlKUyHqq9Jpu1IoVYpxP1WeXBbzRrIooNKsO0kKtjxeXrQ1OUfdsienuY/kSbyWBpKS0HvC
ZEjS85GSDaz6kPTDDWPaSD0vqiyQuqaMQyH9f3VGaWHiSkPywwVZBpPA4itbCD7cJJUatzIw3gZ3
zE+6lppSVJLpTXkLtQfiCeUUCCBfq4oKlppJii9VSfYmME/aju4ZCQXTzKSW5Y8AJuB+u8IQx0xd
xXMkLliqS+NFtR6++80fEHmF1IWpDsD+FLfDeG7A+TsUhQzpL6fg1X+BUvJYdJplAHaXQq69FE4N
hqpvMnGI2bzvQNdSYOLVdgOUt+t9YmtmXTt0gbsxTZrFIMGgc/NLw7gr2XUuznDHT4lEjVjKThk2
CoRubhnwdxn7QBx0zK3s0j6a5FeAY0cqjYnHuuQihIg67cw1B/CNNXPUt3ypyjSH/ZbVQ6fw6wpD
g5Mj6vwzdYTuX9TQynj561n1DFFdEKJKYU1PzqKWlV5YqNLD5hSIh/d9pC2tmNRr6KFskgMWh7yj
cfD+vsbE+seqjSJxOylYSpNDieO+3dSAtbYn343g0fgGOC6VrM2JFfhDJDIppd0dlEiRen8A9/s7
4ISF/yNn7LiFygR8jaxObKZSHQDBN173sTowwMkb5MYzEB1u4pTCrKrcpCDFXqZs3aOhTAjPeV3X
aUqoepihNX3cufUd3Ov5ZbgaKVrySxuh6KmsuD0gd92O3pS6kqYfZkr2kG8yNnJfzY0+8300A8CX
K3y1z4ivmiTZYyiAKkdpDYKaAVprdXYCihL7Sc24Ai0VsMxJOsjQ/jlTxY1TtpVo48rxvmeySN8f
Q2ZjKG2YsZA77xzSzwPFDa6fVEhMCkv3f4SJF1/xEvvcf3sTZelaTz4Oe0IBYJ+3sDYXFgIWzYsl
qvmykMr4mWeAz3v3WyKQ4c/Zlj8DKBrlBgwoUoVu6uKspAmEPhR4IErk88+p4cNvpqOZta5zKqvp
+sebVkxO11QFxGnJkDsQ3OFW4ejdjd8l085R+AxPYR4CqHowzgfK0RvxqjuEuiGM2F9HaweMuvVP
enwD2ijYPnY27sw0UOmhcmj0tN3Va5gHRUwAGSPqlABD0iG/TmcvlznT0hfvJgCW1EWWn0FW5QsC
vPk/6ccEyb0CDLQ/RV2cbr8OVzNtEQK/i4qh11CDkKHunG8Qud1CCNztaVIuRGi64xTxfwMZ6VhY
MDNfoDo3mwZDLwadDYt6sAh4d45UUstPVrqyJK2ZM06IFy/kQMT6eU6KgEEAL5rFiwpH/IVlZHHD
lvU14bUXtqKUpjy5qwkdikMBx4aOoj5dmfcUaoqd6QOw8mhQ3nNNsGQQ69Gqv9aVcSDun4aita0O
8AaTExMCvS+aOgsjbTqkIxsiP7roAMapbuFS6m6cbTqDszfHR8S6YTG4U/GsYBw1YMBMn/9FVaO6
du8PJJYRXESMRPCSedDU9NQBqkQ3BaYKHC88ndbO2gfz+jEppv+vEDWkoCgDqJQ+DHe8aAh/Z4UJ
9uqHYO2wX8/HWYiuqezMiQVkto1Ks52GebLTc4OiHWCgQX3ANemcw/VFIHVSwR8DLvDrsCrE/4c3
gAolJ4oMLtPtRRRjMeR2m9/RbflIfk+mAHj+xitM4b5PmJGJSUcwuNhbZrG7Vus1ELBNhYgyvZAE
NL1QHtD4qGh0UOK8n4k2TOBI50wcVgVEk9vAoex0/t3yaVZ886bQ3oP3W8v0kFA4jVQ1Q+rACviw
DRsjcPdCRRDkrtod0NbOWtSXrPukxs65A8l0+OnBkZK2oSXMf7Kg0JLGHV0Q/Y1Av2i+278oG/z0
eibeAH8OlIawVtM=
`protect end_protected
