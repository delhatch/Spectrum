-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Bcr+A4ebnvpBbS+9KqL9/PbY2nF4YniUtLNxsChIHGmBmXUeBeYYdD9i6p40RMIKZXo8FNpznUkl
X02qi9HbiVcYLKS2g/aimAtXrN3NALKuba9IIH9NS/q8fuSXVBex19J5fznIIWXXcjKAXc9t/15j
7GYn75QStkr/gPkAZto9YT4mhEEcETUQmfRHqP9O+rLbZSB3QpZZcAmqWYK5sRLwNLKYLJylsRz1
Lfi1B7Zr6CsyUE6doXhmJa5b1Q8zQPndER1tYXQ4iwIrjxmzBEWits5tvaOEwBb+ygTnN5J2ElGv
KODTIBcTTbMtlHiPWvlfecN9LZpBDKdhgPmhBg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
QZNAxTBGcNvD5olGx/vWZ/OQWwCldZInTIPcsJAkIEvDCTDzwUE132vh4LDqZaSqnL8tZ5+s2Tcm
NfRMJK1ltr2gliYmtNWmdwmT5cjwmzbqNNfEebILnOEctC2o36L/Ri23FPRM8aMqcIFFZTPVhJ3X
0PdXIXONciZ6kEZTZpvqs2+TTlKMnwzEN8w0iCMxhWzkzLwbxzNjowczqyxHohXWAsj/6EYS6UNi
/mDamucJ3VK5cQZ7j60KySyb0UWLH7Ntw8tq2hvMeLb5O787ibqpGaJDEfPVq0WM5C0AhyXCzcY3
ahpgu8ryfd7vttGkzZee4wmEujMjXqBYoNlQ/kB/gTY49IhnN6mD5WiPKHvK1iL62kQyAFiYjWBa
TOwMO6F9w+ygvQlZxhGD8pvn6mLCH2D4LgOSOFuMlSmLu7b2xK3t86kYG6zBdAAkISaE1FX04PQV
4y7ASlN/nf9BCRg+FkWHCgsbGBl2hSBkLgPg24xo+GTYTcVdbkLtn2k2zQBklZpgVReCec0eOiIp
v4LSuCCV+4dp06B6Spf1YO7kd8bBwvD1PYLJ9rvn+ueKhGeVPuUIwjzswDS8tG1b/3LBSj1ZtPsr
kMXrvyQVXwWOHdcSCesZidZwGh93njoQllUrkKYN6KvGU02jeZDuByXru8X1O4Qdp5R9J40sYXU6
ZdiTcRRpOgX9hXdX3fYflv2h+6XbaF7JHzrEAz7VM2GBtf3u2IhAdM1WepcNw/QwmhZ3rAJxDdbK
23tbEV8D1VWnNQaRcohQyh39jKHEjJPzTG3q/wW6MQtExZEtcLop89oEJcTdEUiIHNQX5w+KRZhA
GZkBCmx0O9FhNARap7R/WecwSC7H750L7ORzIE2KVF5N7uv1zRKfVfWpAszNW/LtSWYQVqt3Zvet
LBJq36cnXIeGtFKbAHSLRv1UJ9BquoJbehixhbcxM1nh50tTJKKvCKg8gqFFmstEN7htpNi+WZXs
NsporBXeOCjbBgBcn4qQJqfLCvV2v+xKwPLdtNuapfUcBIdR48U+q4axjpeDshCR7G0qSdGMAHf9
F2DwPwMV4fDyyH5T50peo1FE+ZVaQGUMNkdT2Qlps5dzTIdj1lQBr1juCF8D4yBVytFJ4oyGB6Ke
qZUWKnVPtVJbuvecFmzLnRUhBFkSjP94NoIVFE/vOjWGVStD+u9tB3VfZJq7uLGMo63D52lDBtE0
kQnxwIUiWg/R1UIZtFaTUXRWdL7FWf+qdlVP4ymiBUHg1wh1nEGYYkZzK35kxiGCc1uwcPsifDjC
JVsxjhcvk7aYHrdfniffxnLpJsK88DsQa79MKsOTt7JVyaYBc3nH56b7gtrsbLydet8kaZgiDpOX
WpM+Gzx+3HN4ldgRi9cSzT01W4DPRFx+219dg8t42DOW8deIfx8zIXs1bRfFo9V9mwMykAUETNDG
pAGXddwutpfIMCgXMhG9baqeKI6iUEma3SF6hedCoi5axWydUoYabHC4lc26zBg0MMF5F/QIvANl
VvJ/VRlLIlkm60wm+uqOsYiU01gnWZ1a4ODmMxedGjUk3ElVj5CNMwpyuaMURqAe9GslOaSnbOFe
W5CFLPgiysgoORMi7LrwEMcmBbA6bRUKCjewWU+QYWrHI+DTouEEZN2Edx9N3EC21kGxXiME5EPu
3q++AaTZMd5uwsoEeUN/NanUgXCDOQHPuIIYiiVGpu9LT9FHndp0CqyD+XvIPBQ+FhfK98FwhBSC
yb4n9DrVKjbd2bw1+3KTmOtX65DGfKK1jddVI1fgSzT9OQ6itSEMAudlSj4R6q/jJO1+4fI1bNE0
I3V8KgrfFQxju/I7Xg92Oh8KGHhdzektEqzLJFhlJI+FZHdjKPxJZ1+n5V7TsDQew8jckuMkzSGw
4ei4cGTYRc0M+HAz83/FFk/ggSpZotfXT7F8rGr5/EWu9lhlPasx2+HtjapamkJtKGSWRfmpbtg4
mGZn51pcDmZT3tZiHi+Bhk0woDT2qVtpUAZ8HorWwEvX/3JdxBtYHZeptoVi736fBTWlqPaSSQH2
WHUNkxGzHpNbDH1VLiYwf2hL/FMzKBDcj2NlATs+jXqO43qGQtFxtKhuLG0yZjtjHXowc5abLJ3k
Pc5je5SYXLuQ6nyf31MlNXzrCpARmkkF1mdu5QjJ5xykXjUe1D62cP2/sJajAHNCfto3QortT4G8
v28RDER1W3K/By/gXKiiNXYlfBtLzn6+9Q/FCu9YmlX47RJw37alUHdDfW0Fivy8bshcMAezZts9
UorITgFoTEEyDKn48+wemyOLQvWTV9tFLgEqrEq03FjJhsKgLyeSYpjQS7lhxftIDhoVS280PGf2
zjvv4nks7R5/kC8DTD9RNWFWizGQW9bneVlOBtpvFPdY10QnaZ6jdhLp0lglXvl1Fk6a7T4uvc+1
r1H8A4r0O0pJ9pNE0ZM6Mv602E7KNfZC/fCLfFODBEMtwOdNEaVf0CWcREiL7v1qdb4QBb1miaIK
iRTE8fjllheXDz9Aw290R3xTn6HzFO7NDAegXNCGJuvVbO+F4UqPBO4AQydSq1wRFAEhofo/jtHl
SGWDMws+FRlHaccNOqGCJss/2CKOP+Rnm3+RAJCPi6mzCZSTTue34db7sXChnkqPzd5MpZ/mho6k
aFtpDiuBBQ9OfLrB1Z9vDjo0/MGmirEBO+cqCn4GGPUbVsDPmIyWtf1cFLPxs3F+LBvvSP6ValCh
wv7FuImJYW3WB6E6n7wAlHRw5+YLSt/h7szfEGO0srjY278aa/igUroFBTXDKudzfXG9Lw1hH8yZ
ZixVzecGqf/d+VTl4tMt1L99rqPJnNJV3u1IQPOlYUzie41+56H/RimwlyRuZAarDml/rMYBoa7R
0u6+YdEuAXuHntV0WNd2Ik2i8cTH3BovTa0UtW0lgjTiylo7rHLMja872G/+geY1SkFMlbCbMXIr
RtfScP/LV/VKTvH+w4aujHwPuEtXHe8ZI5bGg6UJQV6GW7q+jfz8XPkPeGuYXjm2WvwrJECNGEzK
nbIXsFjgkfgfq7pyWzrOL0OHvGrIPeHhU7nw1mQvyV4KDcgOXy7OJ0fzfZ7joUY0M7OEfKgbFyvz
gGDhMnVmXsq9Z8bMg45HPrV6yxugqTX3+HDwZvGCHGCVLU2RJbXkV9yeKxaOjXdCoZZGBiGANZ50
70hMY8pB4cfkEmI+8Yi7zAuwol7xNyFPRkXSYK/vR9u1gjsGXYyrVRizdJtz0EYEhj7SJeMypcqo
DOinKSkC1vRV0QdqjtH2T9bJv8fAC99SeU6dHl4VFp+gs6WCHvSiCFCP3WaNg0UQAIuDHuLYF6iy
safoVdmLdXu/Oy+1VI7/3Y85mfNL4EcmwfuVbFqt1oEaTWvN3yQjovYTGfMfiyB6HbgCh4josdjb
uq7kbV4iR5Pe4F38GiFitSO6B0lyuTTHZY7VAZv+MN5kQeiYL/roc8yV1MoUdOqVfKAxg1HqvI3L
0X/bnOcMjzArByphzuqAKbG4upQMpnnTABJMtpJbsS5O2/bqEm85UoHPSMBXJYjc4MWovv65DGjv
r4eGOAHNqgvcNXU3e9VSbuU/J+PWsT5c5dff74hfqc1f3GC2mSwlZgF1QJ5os2xBCaB3/m6GG5LH
rgNNt237VnbCWblblsITOcW85irtbCd/DEygGsG8GxhxINL/a+gqb8kH0oj8eVSKBfhuxeBhx5Ak
PYERJ2khidN+QHcP7EzLWDdaQ9OznHXAes8JZqtDNaGoJT1GW8zwrkTY59Q6YUwHucEAZp6QuCGi
pb6biUyA+wfNxyqKapbZf3EC5r7gTYkE76RPcOSCJxZl9EA1cfUmwB20i5xRBeLGSytPHEbKkDKI
P9eIh88t9/w68DTYjQIJsDY0NePD3J+mWfY48/VjCtCsMrABIdjRg4trHvjtsVPWjRlqFhLxx9TC
ufyfyqQBeYRQp18Wk7CYSrLA0pOoaZ29A5a4h+hIksaWRn7VjxD6ZBGlowEm+jnViKtDC3nFTJnI
oQYC6Pq8jBtaFKGrv4Lx8aRyw63BbQdxkhXVvF1asyU3QZIs0iM33NtOuFiptU9NGLwizFv0COhF
VmC6Ch4DjgTPNuJJ1+n4TgieZy5zGbAzEfmujE8NCAh7e94ZwGuJtEgeDt1WoyMTS+9IFJPXkx9S
9AZwOax2p3e+nCvW9DX0JJAA9t3QwV8Nazi7dEGqkpzCYlW34WSer88aXD4tzpnu5Q5ZgKE3ceBh
q16Le99jajDjVhXjQM6KgDNyjhOOrKCqhJgSnR8wLBxMbEb3lhSQsQ4IFIRS0E/uEJAWibc0JBD8
nmqP32iXyQ+Mknd7NoBNg6lyUInebgWZBp68Jm9W0LuKZNjp2CVsiH+UpwZcTrrk73UTJKHJuxUU
bCcakG8O2UPnkdDtv1H3OfMuX7ivLEHsAPlvXjqaQ2AhosiBaXZU2Ujkz6Nbl8f1y698MfPwfk+C
voKU0qnO++xLKi8bSAqA4auV0eiyrxKqO52F2d1Qhw9HGXw4EoS7v/j2bxAlTB5bhhQDbWBW1Vh5
YhBBVSaE2Js9kuvV/Tdml+dqsJyt1JTGy0BIe2NhH5+R6DFoNzv6rAQMtC09crIRi7C5fUCBPDaz
UVcYia2j9PU1kzCD3nOuVKpeq2J60UJP3j1yTs718XWiKPdXbaz24R+AZ8Z893ik6Auoz+mAfdRH
70qcXWAXgblFZnso7trKto3Gb42KqgcN+JXpP1Q6LZYjgHvCzun616s59O7Qe+YPz8WntdmFb5jY
MbTUlKH5XbD56IPEjGHZnD4KrJbrhoZXimRoJj3bQrdn8XOHKioKnjc10KxZoMO6nneLoIUyrQKR
uyJJMzpBWBA8q/sZxH2qUPKuYrIg9rAcRiQUZPueR/FjzJMaVO6GPjbxKZBZwqve3K6QPZ8D8HCO
BwqAfa+EzDOiKaQIUSJw+jhGl6Qp/Lfkc2SYM1AJwdtBRa/X8idWu/Nte1kQjTL48Uc+dktT/TQH
yIiHVRfO2sKM1x0wVK1FLSLo/QBIpX58i+PUafP35YosdgvWkMdYvsz6AJtO5/yheuB/Tr4seMQD
v5T5zdZ/FdA8mqGUq/T+d3sYCrOTNJNmM9jcs578IFz+7n8U1M/JU8pZkgxvLU1FtRvZeiERfnqz
A3TdZ5uDibPaWzqUuLGCbeSrNAz/j8w1Vnk1fwtJFHYOurYgtLNqEUTuzHUwZfCx9WKJdCT6avPc
t4CGi8JSGMz0/D/D1b4TedfmQttlN+6SqiB2xgLBhtnMz2OY3oAv0n9nyItjbl9AmMxj0cBxZhsa
eXwun1BMdWXOEaGTx/NAml1BdOMTxvNQIUwcC5u8FaBnLpenxNN9zvthZCPLDBDBVz+9WmBVduMO
MT6tV1SrzsIGsVj2e3n3pFr5F3i1SZP6oBfyICEP6oEVTE1W9GSly16tAxsGEjcNOJpNIi/00pBj
//jdDlsCkEBwJSysQh2K1ndzwPDewAnjGPK/O+nHC2JRjb3VrrpbopeTV+pImBevDNOPXk17urNX
32jdew6UZo+CybMnb9A+grxGhGBBTd9Kzt+0F2flN4KMCPEyOsppEggcWRPrNEypjgmck+Esimhm
iq8jE6p/7QuYlkc7HJoa+hPizGmuoogt5iCCJz9uaTOjrs81tRCq4GjYhLqf49eEVQ7xO1Z3+ZFp
Y3LJ8jlq5D5cc6G9twvWJULoBVApWoI/KkS1qKOLLXJ7fZM4VLdUfdZenx7obO+hcF/XWh6MB+/u
rtUVSAiVH5XLAYnPlJj3LyxpYFQcMHf0oyXNLVVwB4lrBP09fyNtSyC3DP+aL0W+UXvJE/Pjgju7
BDuF/a5hhF0BH4xyzX95Ijlt5X2wzVoaIl0uL1u4rpKUfVzKj7rO2OcOCrmVaISSUBVxIqLBQ8wv
JTPVhOnIM2JhMo89a+DvkEMl0zOwrWmqn6780rxY6BOIFey8Qv67ZutLQY8O7ZRX7vJELHCeBJ+O
UqZTuGRzZiUIC8zmmdX25FbjpZcJozmm1cdToX8cIeNq+E/pFFPvj89ygSDNw7/TmsE8DbmmS5E+
XQs8Ma5O+6LdYrnWDMBTySHnmZEDi0dIcV4J0hbknnqCQxIcjUFgvBY46XBvQz1nlC5JW1ZQWytS
jhqCxGbu7ZBTRTzMdWVtjdxS9G1IkScaN5PDSblsbrkEZCgzSLZbA03wz0VuXejWyZmCd+aG+f9R
YOBEk0OjCrP3Od1/CjZzzeduqWR1LyVHQXjDlwOMw4rFqyl6XO/R+jqR0T2hdjO/o4haB6Zw99oW
AgQc3PohtDFRqTyA4KLhPsk4GbKQoYWVBFlX97hFZp1tePJjvrmX/EogMKEU3D7tpKok8rrcE27q
AR6wIyP1VgJ+kbF/W3+nwHb3YUZcF35WlGyoS9X82D0phapc60BTP2YIajhGgBz3dBGubtyCnWOm
omnP2/wRWUmUL6ImkHDJ0TcdwladTyJL+O/ZoHdclM8ce0nwkt/ht3NJJ+tnnrb8njD8CecZmof8
BsLURfR3pAK9tlbIE4RhyA+WzAYo/LcP/3ZwbFNstMkoIeI+7sZ+pTa+caOLQCaGqELdyLIVXt9U
sc0RRWF55mTgmlNTfdiXVvoZ9BHVwqv5JG1ZKfRjqdHWGUkeCOmM1LPlh4jmItcTMFXIQEzybXGm
PKAi3chB4GOgOa7EzW33N4t/+NYFVPOIo6IBCOL9cofdnyDrIpQm9ZgQLPwpwnT+Bz/1S9ORU7aX
RIjq9zQBZfgKQDc1antUCkoQpGI52ZeT5TavL5w94b6PCmbLlghVfavpzmuxAakdKkvnVtIJ0Xi1
syyy54xdmV/FyVw7qfVYdktd8CuBRLkyz58CZAbiddMh3rp+VTXnL6MsmGhckpQtBuVqEXG/Mu97
KoOCgLt4hwcgXJ4zKtgNBE+N5zMoyO+gqW65mVSzgoqOrfSmtX6LFbaj32zagdJ5+2UTo/WATRPO
m1ZdyVI8CbpZ/sX5fAiBWtHP87PGaBSgd6hdj/LVhHAnxHkF8iQ1LUaLMNkCiS4ru2GQLRWlETd3
1jgZuHKij6me03NA5GDSSk4ZlO1eKbgTqX95ngnLTquiFlurgPbLCNrFBafcJK5apP3illAb8Yr3
AT0tK9r7n/y13/IRzF3hAKr/B7Pw60cs+FyD3yMzj/cfSdaFqUrP5+wa9+DBAxc500hlmDyFYC3+
Fy0RBphJ6BQXZ/D132+Xuh1j8UQjipe/e09od20xqTjmKqHeJISUwZLF70sAPu65P3i6dB9UZxED
zodQhwm50mu4B6QtNqHvGU1hzsVnIGXpjcb7WRSMzk1wnItjNNChk3aG2poYfpG/sYXrCuMNEH2Y
cgtPo1pfz0mUcvkVLjB6SwCrsKBuAdYVoU689F5Gaq2GkhP2fDBdRH3XlgWZKywFMMJq9fVbhO6X
/eYlAvUB3Iw4GPIdsF74P5QpBqtnI4tl1hOtJc8AzuflMqFiEorBoaU0QYEiQuLcCbMDOtQHiT6c
QxnkgSyNj6VBxRS68aX1cZJRt5NUS5hfPfE4oDKWaFhMHaiqHV9w+wjryVztzKD5BjYV0qRTLBDn
dTZGkVOeVW30o+AmjLHp92amsWdEfCJso5FKrQd2+GkeM7YUhKiWrijHHrth6qNvF4Tfx2BVJ/42
PSh59Fq7JeXX5lgqV7tJZhZYOm6u42mLgkiujQtM/Y1BUllGFiUUKOv/9qMHfYj7pdj9JDtDy/ly
wL47M70JPzDHrUpzM+790ABFfHFTV2QmF3PF+wYLQ/KZGwdDCxhyZB78mCB+LULoy6VyizDNQefO
wTWIWhvyDrhutdBY9Zoasp03ZRDk5eYoTGz7ocLvRSoqAvCz0FF91iOMa1ob+CMTWw/i3z/mHdHF
xy8ZE9uHPV827yWt8NTv/EQuhGg3qP//jLwDbmD3gFYfzE2ZePAQAUs8z12KWPJPK5cgRMYfoZLy
6Q6ka/l52jRBbz+6ysnZize7tQG/GWd2YJfWLhjHV4JdzqCha5Bgg0Z/x8DdgnVMf4Mwr31DDqGn
vqvzryfrEs+cNgoA1F9uRI4J413VJK0VodXRSyy45PqxVyqbXcE6cHAfo07P37/p5RKariYGBXT2
feOrEj9t67DhPWy9ueJk9YzITjY4WUO2Paa8quSC9YUVMY0yRJIbobIoHHODb13KYbnbCbXHJ7mn
qzbDyURpepRlWPFkorUE13HXM8pFl351tkF83S6Ta3qbftWWarawBZavZ+1tN+F1H5EjGkeRJVQQ
bKHYlqLl7w4N0IlY1a6n+bAIpQ6bKML0G3aPEzy7zYCY4PJTDoqZgRoBxHjzl5xGSUwMMzrezHtP
b7V3ZRrsGzWsBv2ep+XKFApRtXFzpYl2BmXQQT+YUA/uPVHr45MCAjI5vCWvfexW06IBP7UIG5KE
/m0Jbnj8tBlPvrVw8r22ahltTX63WJ7zmUXK0/sKkd8K+mzXB6YP/oisBvdxVyaCT10XI8oMzLHY
takH8PTmVWfnn0YEw9cx+qZ9kAnwiyEbTEnNPQlKfyuULttWoMl329jDtWy80NEMODs4bt0ul938
vED5tiXma2OntYfE5D7mDSjyTN8sJZuR1re2kHnKDfUfcoKvz9fl0A9PWfR/4Yfo62yqnT30TxBQ
IEZNKIAepeMblHG73FAci/YuqbapJv53+DhsjIYbWszWIIBQu8vH4P1haC0+++IIoHukNxQOHRWf
oNbb+FQm2fWp1HOiVyb0QJ2ptcC1FziuwI9BY8oZmQzBvHrsFqDYBE70pksch7mmSYTQQlxnuoS2
9oWS61LZrYKns390SOqiE6CSzPiq3cMXwi8nRtMnY6LLU9HH8JVg3fUkw1MigV9pFhAijQXIc1ln
YOPaRPJLQwVc4fm96uTWxj63dbs8q82FWR9m844fRfcg0ImvhXua6F+FhP5KTFlEhuQHuPx1Z4UX
8uuh9eN2Yjv6Lb4nC3svAPeU8s75nK4YdqkP2k/xzUaZ3jiNQS32WTMr3+/MPtdhvfOFTk4dMYIY
Kq4USNclRw2fyv/ALZDZvGnjg5sAMoslCenoEbtKdKzd24S8sRv9NldH2ifWkDH54y1Av9c1WzoT
oTZY1lUKWgngPedNXDaEJTOpaAPczdAjuefqOkvGdsI1AczHD4OOLMl7hfY5pyQfY/Qf2ms+76II
JyW+i+RSBjcmvSMuPNxhL9df2wA+LFWn0sKWFTvk7QJacTd1UxzYaldKuNEa7yM66iQZxDGZ0PYX
1K3qo3nw5LmoeQQs2sB18LPBdTJWvDNjuMBp7S6JMZY+Fo3iVh9fw+jdYk/GoXmXh5LLqYMxStq5
Xr0xIcjzYV2nHIDRrtYFFmyt4F6raC2WeZyWRNHi+6t514eQ2AVQylLAcqKbwONslE7/DneJ8Cpw
rLIPAHsq+AgtHXQMqFSNOiV3sSUOkXLokXCWmYgAOBF9NDa1y9oTOsHueMuDfcsuYe7o9pFB36PL
IAMpyKlIBDPL0i/PKBNTuRbL4MjjkVsTzpyaJP4/QmeD7NH2BTdqQg8XhDwpPFwZkQy/dopKZDE/
m91eleTaVfwEHnFuMjvpu0RQarnoYqkMliQ7khsZXWkmqGDNM4I7NuBr3cjqSLPcM1etSo+SpvDq
41qE+K/vkOsIj8dBl+t7Q8FRVpAlfipt9Y20dky7+EeBUC86lx+Cc1k5ypHkk0olxCh5qhPy1kzz
m49Ybjv32CB1yqaz4lpo7t6P9StD3Lwbd6hH2sjI78V3i/VY7ENK+2prBJRMYNhQgsIB1Z+jHsPw
JdPAJKo2fAAYsxM2Ul4iUFXB2voVI6lWZYPHPgEtnAEZBtLUEhvk4P/snuJoHXUB6IgR+RCJ23k+
g2OR6R/rePd3+SHvCkIrX4PPdW4m2fTLSqHQEFc4IUO7DR+Kzln230khqHB4jC/K+DiEypXB2nrl
dVX7D0UOJiHsbYMAWqRQYOqEs4T5qMY6FLSAIa03aMGC5X/ZtKCxTRcN2BuoGxOrBchoaUGXsEUv
eDoJnn0HHyA42evYmZJi8yeBf7F7kgg+1USEsA+iLaWPK9yh+k3IcEYoh4iGYagWrcf8Es5seRik
1jsigIExKH4gd8/F84XZbBPSAWryr1Fq92f6FQzL13j44Ot3DEorz2zFSDbDuISSIEFc88qWDHq9
u0BmsNDVPS66phhEy+qHCPACnU7Z5dW0cQiWNbSs97iFoosx/ZmURCee7J4plhutgphFtzMjj0Ki
a5h++12CWp8eg/7ZYWp7LwlQlY+s4KMKiMs+yjyj6KA4Pk3vf4fpp759bcWJMJoKiCOFIALt85w7
oPveiuEa45TaO4Xea9pQK4pxCoMryc1J6BVJTRAXL4p/lGYEsVZAZz5pOV7/9/T4hSsWUEn5Ws05
ez3Rpb6+5VyI2z7HpB9ggS4RzJDB1A0UVFnAfEhE/09Ob/eshHZnJPQK9wXiStTLUhqUFTj4Ffat
k6G1kzg7wcBKEeXErdZTeLEU+TacKj/H/5KfMogUUB88SGxMKv8rlgRWE187uQxfpDmOteDia/tB
ZjFVCIA+IskaZGWCCQGVokY58rmg8KBZ/PT6dQ27BUUOEhHeym867uCcZankPo8hESk4NBzIr4zG
qJRxUfbjDYRUUR56PpelRXprJSINrQGVOIsRdFgUJt4CWz2812KYDo/WTWH85+ohx1g94lb2aSGC
U3M24bNneRQ7rRaiXVWqLUALfYkZeb+KSZXZJzlrOv7T2dunGCvrZTAmoOoIQlGNCRdBiHg/KWzw
hvGzuAG+6KAQud1fbSSd1a3xYExXzn05ASdh2xXSOOWffiIYP+c2n5/jz7oALTkvqtJhu5UxVIPa
/S8kFSe3W2PlyT5GgRa8AS3MVmWogOLOe81L3LPXIe0vwtVyDIS4imxxLOMa49zHhxAIYVJfz1g5
zB3qhPuQDl/9CDs7dQyhOl5fj1z3q4TwiuhfhSG9FjEQANdMHtT+ooyT2k5yLi5zLh+y8/fWD1KT
no+cO3/mZCTqqNzQa1xmF5RqhYk84LU8o0S1IgzsRsUGambFrqekgRYIpvMtHOhy2d23EuIIC6Uu
9HKpdObHlHKAWYlLkgefcEVQ2JQ52j0URwU+d5W9kdkORxcfeElf2enbz21QvvCNvV2RjxpfRfn8
oEuKkknR6YYcRbYoYdwejrxupHM4Ix/4dgd4ExmgPUT7+3qYPbAFbpmoUKWQKnwU08r41syV2/dm
lmiwpEqnDmQHwmrFasQvcc4oggaMgJADdlwsUUI1PEiZxq3Z4hWe8Z6xOqIx6IqdP+KfHxpsY21n
nvOFEHUeqKxxXNvWY+p4FqJo3PyEOLVJ9g2p+sAY0TfSP7T7VZVmTvujedt6J+p8Nl0Zy7nGezwi
RzvFIYn5G/+TAPay86tYgBDABHe7yvKslG7FaRLaUhKCOv00ap+K2bDrKJR5N4MuWD5VxqYdZBr8
5ZflgkmWzKBTUG9BdBdBtM7Ljgy1MsqhAlIb13iDQ7qqodROXJLFp6SU7CVIrbf8mkvxo8m/k3PH
mannw2Z7ugPCzmfBu4DRwxh6BBbOukUfZnjYTbaCplKpjsgMZM1VBoGKlRapvu42edwHb+RNTSS2
cuJmvcxP5BMFrW4SRAqDrqmjslP9QRZYEV+07gD3Q0T6RqtIkCMQo/3It7umvQsPusG738Qkt3vD
zYXMWaWsgTvuYzNB1d19kdyOanoG5Cm2jBN+wN194hYnfB8U9ByPOvxFDrVfLgiUB1CURIgKe2y4
tZvj/QU1BVdb6QOqa63L/gnWhXxxsQ/8Q20dGQ9FqVEp+4AklQnWyFehrGsjGQGVlGF+RrHkRDfp
T6pPE4bJcvLvgZx04NgPJEh2hQgecoyp6d+zxCVVXIZyfHxzkz2wzjRZ9PAvsKvQSQz2vvMXl1ln
ecF41K6FdGUIy3UQkElrGvq5dKgLzMJmxz7utNXgPoCTqHQgoF1qr+UKudY9GmIROpmb8DHQVvPf
ChSdmt1vHrt/VgNhWQG3qTeDzoprtq9klf95Jp7EwFHSusMM9XuRU81H96MmKdPJG2CkU6T9/Hjt
H2wH518vcKHeOtoG3pc1LVe6IX29YVa18/O/E0kWUhfTwG7D3h5NS6lv3mgsXnbSBKV40f0b2qka
9U80n8+oFSElrM+mGk3BBk5Le26SwfDt3TqvwbxAfoKdWwH7CnIy2K29uv/S2lQf+vgQyN5jW7uq
0sw0pdObjvqUHj4m2qn0vJeuhL/30uShrdB3DqBgo91+X3j/cKAQ/y69yKIDbPazv5iXPYLad95v
aQNvtzqihGq0MIk8jFurwF6Jl5MFKMBVdlN0MhoIlHTIDcOYB416WGjOBZhnB1JvsGDydfT90oW+
yf/fh2LmPqnJua8SDGeEhTQM088mS23cLK9qf3KOZhspuYtvKKmkq3EhHzvuA/94laCazlvVO/u6
qHFC0S3Xof2AWBM0rYZ/0yndYug47d4gE7sArKStUw1+0/D4sdtI5vNzTEDGerFd7YqqyRgrxTAV
PT5hvqPv0dRgWsapvoeREnMP5Gh6MWMGawbd5yA9HlSKcg94qtBw1r/LTuWophFkLR710bNg0o1C
q2r5j8bEaNnIZMAf2oA//k0IqQMpFYwdYXbMaMep4L6MRtdfjTkR7GwSlqqk9Rtq98Vwtn3TMhAT
HRbcB/zPs9O3XHMH8HCkmLPURf93XminEvRy1jA4HJw0f4GJu6PskgzmKi9ZM8xrRU5Jj+8FXHKI
gd1rmsn2fFGbvF0PIsfktIonpz44MFALu5yUDKdnY1bosUJ6NrHrzx607Cb0sZg3f1wFHAFqsvUS
Ph/0JBKfsCwFd58uUFhZL7Kbgsi+WnGISxN7XYexeFP4Jt4AWdq9Xd7CLl36O5CfYnik1P6HEDpO
PEwlvg7fMhPuvtqTrWdCyCeAC3DNwluHRMqvRJGrUVCs6v0fvH3hBVa8p5kasuSqM8nfkglOrMaJ
5INp3Nq5nAjkxzVJquunC1TlwevFGqb3dXvo9W92z96VKpHpcR8y7lCYQf4jo4PEebKtXYiNDKv5
RJSjl1Qc3yo314vGSqFtDgyD8eIQsc3U5C+QiwJ0SVjHKoHipG60S0iQRiySfbWbwdMAFIdn6J7o
kceJGl806ajypjTwvsvxcrQKILKpJOGQlUqORRIeEkcXNY+WVOty3oSmiffYeMwTU3YmN3isDf0E
Qv5qi/e4+1n8L7jSjL/WKtAvMSz5LVzU5tj92F8zZUi6m4CZL5/lXUBNgfSVIaK2VLokRCaYBdiA
kHjXx8dplowla34R7StQRttCBBKffHGJEnQq4yZBAm7b+1gc7Lj2wvnoFyVeEGHaikwHcEMt2dTi
iAMPM0AAH/cRVhytGeZFGEE+RdRZzvmerh3OPAYcATuyCLJELvt04gul8E69ve+WsCO1FcsyL1zp
Jke6DzYrpuWjJ5Lwf35Vtgk1E3zCJ9AOWIdLusIAE1gE4AoKWUNlnffnI4wI1/pBR+KxH5PT5bAN
eXrb1D609LexhDwYbhokzn7xMIZSXvp/ddhKVHZWh7jXAp6uhrMO7d9y3EQr6EIZnpOMqTSnbwaR
G7QwHZm3ulGyjyFRwDAwoO3YjeZiibSQnlcuuOM7AnDghs5hTXOn8R2UzCjnxAEdt7t+pSrOwGgw
PnYj1pKQCCR3u1yCZM7LQNL1jw2xH4ZKvJ4iSqmwIUTQpCTKrpbXDVVAKBvDwAyM3/iiYADlx3Aw
AQRSt5U04RYydC8v828AjShU1pFgNiHVi+3y2JvN005mUGk+nrEkbSIZ4WZfMJPGhrdvnlrfbxXB
1LQyszc4xFpQlLKsJKQoyWEN3FX1ZLPo7n5k4OT66QYFukhPpKnSh85OrZkxYxbKQ+ahSPvVh4XS
1tSEzOAoI5h8s7FpaxLx1hCUedG69twktAuC8XIqgHEdlqAsXGzPOWueFjg5YCMVnppI7U7vELyr
DPO9YCXuCEhbiNDfbwRXYbb5UEv8S/F+z+7EdF32hVBKSddy3jaZoVaB+ywzvZw3QZNVWIHU4nKz
/MUYL44Vqj9a0VDrp6G+gBjCLgZDtjjo8s+7iu1jFHoShNSSm84h0HfxoMW50apiq/snUYUSS+ZP
cGrAZSPrdb25RsBEcq4ZCdVi3SsUCZH+46roGowkhtWqfnrlbDGshF2pIA5Cao3l8mUyqP3ZvTQu
zSVVYc/Q3sdTmp3Uxk/kKXUia9wbHZoJCCNv6aRoTVfQz08YUIt9ZCNSG+TDb64sWSc5Wo56vSp7
WtMAew9tn5M1F4aWCHKV4e6eewWg01BmVMG+1rLVFXAkzc8Ep/gG8oHRW5clOjaaSl8huHUCYYRb
PfNUzZj3lH7xi8frZhVoIy1euyX6A9yjh8pywmduq7tCLuNm1Ua73euKeXxkwMyc3cNeLke93U+O
p0B1jlRxcBwkjm0414sB4xGaS/CLFNUwjTb7Zbh0zDYA0EuWP1fChCmFUMGyft2BTjpfrxn7yIFn
QD1s67iusff+RDOG4fc2TutLxyrWSonvI9axJIFtMMPctOjFPfI+qAPezmvKKCvOCPOCkvVqccuD
HE/w0Yyrq9DuVpYR9XVrEA2zwORfovjXOMfEDepHwHKqCMC+kvAz4vC9t1kRZobtBlYgPSEI6UBa
ILoHfrsQeLR99Ucl15qB+Fn4cT1e3RzahkuYYUQNcM5aVo5ELC6XrKw+tk+GjbJWzeOFu8O4H41X
RvjG9uLHOjj+snMwFUUD+3sp4ycI0WMpuDm7Y6A/l/GXIoQWqwC31ddRI7DBYdV+AWklXQkdW/s1
cN36TgvATykh2HYRaERgCEuFo4yNh1xSGBUPkXY51UK+tVzwJuNEjagxFyfxuryipz5zYYAeUtJ/
1Ah/JG0q9iF0MjHF1TeTxTxqD/bIay+wJoZEuk36IsnUTqY7EfbRHu+HV9mBSc3nBjr8R/3Xro9s
GdNw79a4Ix+KFgi2W6PqTj0WDIlyttT8Ix95mgtmoPLNts334AZX0qGSXVj20rYDGzhLEI4ig/4j
aB/L+DsmeFm7LE2EdEm1aa+xE5mkQ1sZoWUt5oaoyRrN8evzxXNbAdJpp3NYI1yctiKExES3ecYQ
cU6UnpAbREnIjD9ASlwE15uuoqysZCUaD45CAICDzAiiItmjNiHKtpl841njsNsnucXBBBIez0vE
eSstvcapqWbQ26T0j2CGGdps4Op6NSiE6bmMnYG/ddHb1MhnU8vNWO3JCUQCjKn1wziEZAyo/yFw
moVcYWdfSlFQ5/J5pWW4nWckC/VqrT+1yxjf1r/i7sOPS07Et1hPOx5+2L6W3soj4HM0rIZBuQos
adrCnBnz7tKIhYRvbVi+7uCBAwMFgtq0pLF9xOnzSsTFofMSkUvwI7yjCaQoByT4nyXoU4h6y4jx
N4SoiTlBsgS171glZ3vOyU0IFYoJBsnK0TIedTUccSv/kJhIu8VAp82BgWGi/veXOiMMmqL2gLW8
RycXfhVGIM+h/7vGGkjEqqYjwUY/JTCT/SboD1l/O5lkIhn2nGsMGx5ttFxBcSkt2QuqH2a2/CyZ
aiZpFwInhDKJ9dLZJAjcaGml0gWootrG0SSQjHd1aO0owoK9c/pWlKFwrDv/BjPriLkCVjNBb/YK
T17I7tBVdq5Zb3ld+l5HDLlmGXvqbWAeEk46brM37DdnQ/VxPvRcX9zcRGTs+1lOyeSYDwQzbQEj
YBScIP4lAmH7hxHvQRuMzLXqsKyPT8I9Kryyts62+6r+0n871F6+5tnD7qNjg/ZyZcab3xgxuR36
xieV/rPUYaqDib2pM6JJy5vlbGol0HO9wpu3KtZDnGcIjoXmH0CgzI2Z6VDSoOrr+xufr2P1Jo6U
38cklrgsimYLfZc5RxoVdLU5zQdWeUdnE2zJbcwfoD1abF9/MZqCcBFLCiqpNjAEdiduHOcDju67
mVWOFUPaoE7Y1z7m3tzMCql1HuLfpXy+qL66QtV2908ooH9zCZPk97wMBtgQ4swROb32PVFBsXA6
gB3/Ya5ORZXxxjZ95tRXD0SMv67zwFH8xY7exFWA3Xhc5qHtO3mld+erqsFl7pHprlhMCIDr8FLY
szfQh4/9FkbfN+A4njSdhBUAhIKVv+plQ63bYAOOoPAv8PMSsfPA3bGZWsOq1qkj4tYnZjXq1yCk
83w2s/QrGioBQTqUrpEmSpMuJ0eEJ7o2cPp3wsDnwv68XaKCJFfOcMCoihIUywC52FZzPO2iCew+
vqoFM7ScBAAgKl+tHIewifKXWj38ZV/dxpmHz4oUhSuYUM7Jm+a1Sj2XhrPb3GpW4K1Kad7TBnyL
svLELRZ8bYHhsFVvU2KYV49K2DqqRnC2uGn1Ls53wtMFZ7vLc4xYxBJ3e/nOYAB5wbiK10AgzczP
cqnImFMvRufAKwZivms2wMKBWKfU7Oj2NqcXEKn5EFT2TB2lCcMlST83YWDZPyhr+GVLlROJacZ8
ncxgI3hFbmQeTjK3xuyVxHMKf3Z03Q0DIP5LOFav8YBAMsC0WOyaYZft9pRj/bxgig0YAguvGChh
Lqi+umIRESEvRwsISBAY2j2cT9uzUsl8au8QG388qzC76d13UxwrVB+a0/eHrcNQnglnUK8sjDXV
DpBLwPs7MLuUKpbYu5SiXuZeegWHjipZQqwxiq3VYAoBo/vGHWM7ZuWMPYz5bi9N2jBCzibTEzXf
gaf1igClbPbqoF73pjAQ4xq+BC9Sk1KVD22VdYMaE8dqjUpLGlkSAz71HoolX1V8cgwCJ1zYsBZC
kI8fR0KR95zAtpuGSpay3POf5gRksFU5lsmsE47ZOCZUB54TGE+Wc0W00cZRLaT+DygJyoPvnhrp
qq8D45Fy/StgQDvz5IoL1GUesdXINCOYw2tczAgE0Gq+oIYyVaIOyd7owrPbYhUdRpG+zaez0ECO
AsckjG2uxkZ87y/3YC18TkKlx4uKtJS7rnVKdu1TzLEqzuRxfjCBK4y6w7MjI4qSVP32z/j6g74i
k5KESqmYs+wQ9ycomLpEf1ZPJnLeJXT2FttQfJI+58b2nO2PSRoqw5XarzFNsqHl2+spLlbPS3Ee
Lyl1JK79DfeEBPSsfIixQuHxUCRQCdVpGo0iT5TtNAsi6cskcrevZZvdr4Naed6qt99Hngww+KS+
NLDbJiFIxh5J2SrVHCu2Y56qHTCnNj3jSXiuCP+xB+QjwB5jG6JvpoilRNX1sFBzwea/UqghzEnl
fm6JLx7XaZ4gbkJeAADOyvOdOXFH1HlR9+hUaIPQqkRO6MoPGvlUYv+rANYBf4Vpfd+ZfrWLHKI0
FsDz+hEltRSmXqJ/gjESV3Bt1vbx8HB7Mv7d1DA1hjrvepBc40moaFAKgm36Gfx5eoH9lLWqphn9
3H2u403SqvCf39FsBQ5pA2zlcjFk2kl82ZmeGK9vgf14F5EEmSvd5XjtT5wbKyCWwSpDf1gcyd6n
JOG25o6n1u6j1N62J2+g7hzmVHkbPelf/J2T+PblOuZHKTbUoHib3dTz2O3sVe8/z+IADpDe+rxE
3rwTeYZtQVbeoVlbzxSXak7GfR35QtmEo31Ea13D9X40xsTmevCgAC0L2HDtfAhBL80+DlKknzJ6
G9EZ3Ow8x9Etr2ErYy/BW/XzUIAm26LrzS+3nrKkObg4i5C+RiC/win2SsXFwZ63I3JzRWMv3OS6
FgP+Ey0rvBuIbpJYLfga+WA5gxMuSQGLKE3RoMUDSAsdFrCl2F+kZ3Sd7nZnCL7tiQq2tvir65Wc
oBRvdOztDpe4hQTpZ1PGDvi21RzHGTwfYnciNycf0IhRULl7epxe2KwPt3REh3NIsAiPCtKvZDcV
WhnAdSX00MXH0UVc1eNONZ1JTX+/yYWtWq9h27mngwwTw0xRj/UbVCZ3EPvqssUzPmT9JT9xpdrN
6Uk0XyEkFiNrV6Ui0YyBFkIYA2WitsWbcTvROemdPvXZf05+uX+9ANTIZsjLHQ6lYRQbnUV+Q33R
woUb/g5+25ecsn9rOT3J51p9/wL5MJTashVozA2iO2tUXey8atWvpzRrJeGdKSA/13nyEXD08AvN
G+ZQQyC3C1foiU1p6ZeQJKKq8TPmDgDrINtEOmmSbBiClzuyMAYnq54cjZRbuoMhUuLyi32st7kR
4cbvtBKYSw22b0xzcZKaBq1alfof1f7DxIhziha4Toj5tnIm53QdHg7Xq6vonprhWC+VSusUB/AF
nwPw4ERXIYlFrfQlzx8v7Rsw8x9jTHpR9YJ07i0bEOkw1l3bBRyCS8qSxUvIQcMhTh/PgwGFxKv9
I6UfC8c+R+RJIpKtcFi1syepEJqZdBqds7unHLB6fuQdCmGvEXHrcqsELSiGlcaEMk5UpL7j3AqR
hKVzmX0qm8zJfw4PkyHbdhSJhZgAtW7xYPNZ/l++I07n60DnioqIiiER9CsnrdsRJB7Q+e3BTcUO
bcB4x2/2Gj5KrfHJZSLbCuKeDy0T9sfrWi+j10Zx4//tVeirM7dOgV/J7ZVLdflf9UWqUC1+SL/g
FdIuL3UxLbzzAEgYoQ7j+xoqHGtTLNGIP53p2U3VMNmicKGikdbG/4fdgXItBXQnkHNkwAAsmnKV
LLlC2C8NeuKuLfVC8cBWtWKZFFoVHgiX2vPszy4ck5iAnatL3bd7ECwWa+2k22N7zkkKM4dVpHT1
9j+HZNQPcOqV3M6A5Uf7FWwQjhPQIHDzAQ7GnQUx1J9m59j2JMbCO9YfMNsgsjcf/NxuU/tXuHD0
8dHX/wwnrs1Rt9GH7yoqJ2HyPjSLuXJW/u7YIu2InS33b0boa4VgRJgYFZBa9yMIMZpKTpiwSWIG
sDIHGjhBWMCwOkI8lOTBY1bqsuC+TQ5nsXa6iFLF0WTPBLSlpweZFdH+FewIL3S20Ot1Cm3ZgIN7
8z3CNbdB0UjoRvc9Dvh4iVvXT+gEuHn8UsZEW53Qv4VxaQnb+dGP2RM2QcjJVYkYBjmGMtMxX1gb
j+rrGf8vgjRAXZkwL6wBvWJeWOhxeNRuPhe51XN+5ZbF49hTzH3LvThNkIQvKjGk6FP3zcKSB8KO
jMpo9dJ39Zde6RmU683EolnzOV+iqJuTNT7DynfCDTXXruMZ8tss1ncRBux+/U5cMKqWi4Wga1ZA
K/FLYmvhbL9ilWp9ZqUbSpiXfIZx/Pj6vT+GvEI/lfCu3VAsrd5E5jNE2saXfTf0YGdTE0nQ2hy1
BBy8hfGPxQFLviLfkMv1i0qIZb2F/bKBgCwEdQamFr0g86FmHPDP93Fp3jKQ0ia2JmDR2NzhUuuK
a5bkl/jJc8zTEmgi1MuQw7t/pyKGzSg6ZspvVxFfNp60XYfJmUZZ/lkIwELPYm0eK4KrVWak3bPo
WyGnTDC2IRSg+l+eSMQY1PZUhvVlKNWbCsfwQkkHbAOVm7M09dzhueacAKRemcOui94ZrnCSrOoO
qd0OLiR8CZHIE5hdrQ1PXR+x9O0v39+1LTH7h3C0Mv1IoGAgZRTnFq48ECKKGzUHFefcC4nhGVvI
TvBuJxpysbjW7zL2cVm6K3omNaF9l4Pdr/cDGBhI6NKST+WvjUOjvWvdsNIr6SOAvYJBgzhDgkR6
x8peTFr1Bq5k7tRLzRPVlahNNWGe1Kpsa41YZ4l+PuVH+HH8oNgcNV4NbklURUYeBlPLQQ4zEolv
Ak5jGV7xA4ZTSfLTX9KqzozILzdgwvItUmdf8gEY6f4WqtiC4mUH2tVjfJrBP27ql2vYfrdW1MDq
nPPHBa5mhi3QMSit3eDcztDJUSgT/tlhUM9XpPGRVo4B33ffmFMTEp1fMd3biA/U8pXLE/LkuBIy
jPUkOgXHxleWLaKEfq4OenrRNpumZl3gRbzZLjquvifDVB/0sgsm/yOv4wh1BhLCdmud8eLDtBch
eNybmrUbnAMQVnn8WJR+rk8vd/0p88rK5+6NE+J0xNRoqj6LPMLS4IjWgUP4GOnrwPtaJCqVGDWG
irlHxkACUaoICSPRsyaaNZAKjl+e2HjNYLQzjrXcj1dUOM+3Okp+hEBIBGLorONVNgi7UOzu44LT
hX0K0snUokrDpqTbTmu1+XJYHarhDKjD2ZQKY1ltKHVDRUc4BUroa7dOMJwda0jPGItORNlklot+
Ot0zvc+PS1xclkntht4DsxVQE9KmuqBnNFa2KLtr/3uWGB7a12/7ECPvQRCViLVSQCP6kv3+aMQ4
mYgNV8V84a9gVzTu0NgZR6bAxZa4XCJl6lwCPjrYotA09G2aFOTN4yoG6ZkpsANLkBPO1OrAlGb5
EjbURhr+GHTJEkg3oXG2mahGr7gFokui2gZve+F7PGzGi0DiWnrHW2twzg5+ZPt21SawnPPZ1WWP
XCvNY7y2cjSpvxPM1TyKxdikaSbQl7GpuBQN42VvchaFmhIFry6TZQ0UwE8Cx/q5Vw7KhNf5fzOY
kAf9CdhEnHQGtzaPDBXwwR5Lka86349QGMs3fJVmkMAdcfIGO4GgqxaB+jlPk0QzK38z6pl0voHR
6fXG8q5hLUNc3GAmYAt/FQxj6+RLqmN0qd6Lp90NlunjcJDtjTOJ/+iUNa4cdjqsiiL2vWkfj16S
eC4QhnF6xeNIc3jjS7zBKGdRulvJk65CU259kvHg5rBcUX+1ayuQFO3oU9kd+Oc8qXZTgwXWqrNx
LJcdfZKLQC9n6LNl5lp707KQqJUVpWdcx1LAKNmvoYkS6eoVDQS96e612V9sZ712d1KIjkuKROzI
M4JAg9TlkuMG4ITXSLvrx0r0BC7LhwiHqnKr4SqQv6cCUNnAXGH+Fn0N0D2idXT+trQKSzpczHCK
gkWP5VZBrUpGUL0A0GG9ozo+47OvJTIizPtMN37Vn30JTb72kh10pdxTAA7Yl00VW/m1LAwXbXDZ
R91rZfRoqcJ3rJyrLTIW50j+5WILOYaFwHpW074IW5KaYH482Ywugr2yUkdifbdTIRdiUR1wQRNJ
fAqxA2lsAovf4Qg0L4XYI3m3TJKTbyA4whthq67w26pM5ahSpNC8Ccck9EEUCWXIV81WkEz+VEoJ
2gsiFp1r/Hp4yfqIwQieZqyQBw7LPRLp+oMICgshYnEK88KuokC9erzzObaVYDmdJUBGAzYWUIgE
WMnRdQ8lalFaQOaBZWa6WUr4cSZU5VLSdUCeAyztPL5DkZ0NtVwq4fxfc6CA63TFdcycc9mefwNO
cPosJ9O7MUfTWBf7pQc/8zc7h/Rh1bLqiFiHTil8/3vZpbm8dGRi+P2NYiOy0xcmVf/+lci/IxOW
NSQAPQB4cnG3znW0njsRkysYdaQEswivDxCLvR6pPXYQr3uoK4XN/Ao9OwXxUFSS0LrfPCCYwj+0
a4NBQNHq5IUM15DMyUEmYWFcZOXnxObFVgV6WQqtLNE0TY+XbRNUqEmSchn6hRcabV9i6nKvJUF0
33S2INfsoQHGjYr1QdygV9/kp5blAZUeB6Nv/Xs1Uu6y2ghMviUXzOU8QBK3meUlB3Y9T8TaTseD
Dd/liXBkvWfD6sMspbRMMWiqPsAz2XM40o7RJgOD9uo/jiQQyAz6vaC0/rOWYYeORhSSXwukPP3S
VqOwyzI/5XPoO9AsPC0IHGAcixeLebimV7cAFREjumKcWd74R+u1rK4csf7ZAs5kXTzYvEAYa2MS
u8bBkSuBq55Drpg62qTOiLyt7qAet8PfQLV1nebV1/ze0W3a93EanNa2yzqbJyrrGO8E1gYFZt7Y
fzuwJGq7zECjmmDftSiZ79LK4DG+N3IS7IpSIFiHTW2XjKjxIgDzIEBOPuZcSc1PbvSAAPh61KKx
HpY8Q6hcSKcD1zFN+H5aYBtR3127P6w4AT53oxkY0MlH9IUbapDKTPogUoR50ln0AfJ/7Qf86qqw
e4EIXhRRi4bn5KXGhm5ycXwVcf3B4k6/0qINszdc2tsJjEI6uBHImSD8JqbpNrCEtGIcscDxNehW
FJlhjeOrOoAijuI81q0nfpyZA3F8Bt51X3Hwuq5+wt9lZdYxenBknt4M2RYReogu8X9tcVwl9FVq
m5V3kkKIRu0jqr/qJIGi3G6/Q5v88uJsr5MIpMyc0VpyKHBlyvirDAhm69DBz2k+5+d4Qc5oOf+0
EFAyv8zGODXJRtXPm1m+Pdvjb6L8BCGSejKZJTgATkWWR1pEKzwGYMtDZ0FzM3OOSjbH7WwNOsX7
+dfXjXFn/EQNkm+Nw7r3tl5dNwfIepbNNcL4PQF3I3Qi2j2FQxrDrqJhSD8bXnuRsSkR5PrjypFY
RY/FpJ7nYP3qD78A6vviLYIPsinJHCX2L8d4aXXxVPQ3aPgaTjh+r9hGRhacDtgrUTdKOcrL20S5
jGTJuuBE7bF2Lfd7mA6wcksWj+f5swa6D7V7LWtB8lOlazw4j7mWsuAygCaZgu8yGa515aMHLoy6
R0Cw/y/a3G9WDntJVubfHOD0jJuYeqGwy2Wqmzic3H80NSYwbxqoGIWHF1WLT1ZRfxGcp+ZcjbY/
W+k8VcR0Vo6IJ2855jt2b721ZvHzKyyRVQco+v5oWZz+4YK60CQzJQC309teHmx5+/YBDRIHngLn
C81LAnheMQrxCmBRtxF6mYzi20EXAL0X+vG0DKhpHNA+8SxzEGk+T9jCEm12BdmOS0stbhW856rW
eoXPrFt8L2JV5uzf3kFkvkiSvmEmZ4LPTcHVQfb7kvBAqnztc9egO/GPiRQ4GyjnNfDoM6W2tYE7
pjOQEtle0LbS6l+baE1/i19aZJAAo0rNVN8kgyflASQ0Azr6ZqK0KuFUP8m5T1oz4/Ch08/3kXFf
InZpdvobOF9nI4jejLaVcnaNAbWwUT9RGge2Gm0HJIRjtzwR+Q6YJvUvK3HcfV41dIzf2Sy12kzO
QLFCYoC/bCvSeh+1hva1DEjXv/Z4qT480iEo63VRqL52muIz7l5vYqxp+Lvv8slJ3E4OVbVF0WxN
uF5+51l6JJ7JGpzkAUoZN8585bKhfwT5JPyA0wWkcC+s7eX8DnuaWK5yuEfcxO3fHPNNAJPuHrJJ
95ylM4Ju+6++x9SG635j+wEE5iKpeMBXNKELMYy19oYMqv7W5zBZWdswhPkjrG23O+eitDOqJwK8
sbqFGrJWX2ciK9oKAKLRh9hTGP5101YOBIzBMFL8r9S1a2fJr6iuXICRnIcubLf7Rw8WN3W4nv7z
ljtrvXwA0OZXsOFFchfFM8azmNAP4Xlaz79NorheLHs5enKhYOw7JhQI81qDY12PlHWklfFcSqJp
8F2pi7FJLHctd7Kqjr/wcqsKo6ZMqciJ3bL9e9lFRDp+mw46Vy/iRQg9t806fOVU0nQAHnrbHaUR
HumhvmuQv/bjHZtS/sBj+27kZC3zXc2nUdU7faAa5/jzMmM58U0gYTcB+/bGfpxXA2Z5OpS5FEZI
obh6Ki1/BlknLmc84mSsiE1T/Nw6MawcBjvETvCa8anrZZtiJ6KRV2NrDI0kxMN/fZ4bMnPkVnh/
NHqLO+ky7Wjrx/MWDzmLBYfnvhLzxXm3mDp7rl7D9UsZ2zrVrEwOtf8sknFkCrLgHjxwAcAWaEoM
NiKpNJVAUQj1fp2pFbw6sTB1/kgavusGWc2mWrNPQZpPb2Zs8tK5Jw+9DdKdhy9Cac4rt6kzTKu6
0AU1BVkhcm+ge/JSl0KEtXLX6VR2JjfNFHQRjxuJEvmW+/yKdltYB+EWjDtr7f6hgSDecUbttysT
IJCB2HQXQ72l9Iy97ZTaz42h9ekdKQqP3F/4XZTQJ8CB/nRYnRjN7RiRPC1AKCun8xnqrTqEVZ3D
EVeJ1PbNIUlyR75pkzZ5xBaTu9A9+tsEKyCatTx5Jf7Slno4YO08gBYD770C9U95/NaCiH2gYMWy
3fH1ZEfmzcWW9Iik2icUxtDELinfCJy/1uGq3vW8xGf6wd1LhfRkmu3qmD0Wb1/ImpsvyV9o6Eox
hok0FEDgJIIAnq/dct5XwadTsg/Cu8Tl8ZYJ4KD309FnhRbXUDu/RHu/SBmRHjsl0csi7C2pIjUl
BJGDoaUQyFERxmkxj/PWihH84cOJkmeQyJKOuxo9N/F/q/INdFmHChvvfl8E5LufGswDOxAPKv66
CThS0SQ+KPTkSWMiLkKd2WE3qx/3oQ6z9d4PZlhuP45uCVfe+HiXkSOstBlfnxJTXuDH42RcaaTM
heSemFMB0qUfRhGquPEMeowntcQXr3LTq4/VUfReBgtx8P0MUe5i4r/uAlUm20khBYdLQRfgTZHZ
eCqYoth/n1/yRhED6puy3xOOth9y1Clak07WyhwAg+vmRRtbIXvSTGl8benJqCNvctM1Djypy+rE
dR8aBL7pKUp9qxFOG7dyYDND0hJvS/LcKK3XSmWsN5oTf4Jc8w4ccOEamYlnX9ZEU6EqQmM2aJrN
gHbGF/Y4o902SU39Kyy6RdLTH0AmOFgs19XHvrxz7PEOaoMlMausXFUWkTuFxIz9y3TE5IbiyIxj
uW9eWQNFXbY7HaovBlQjDMXZ26KsSRF+Vlb4MVCU0fF12tolnq6MSGXZrxW/2ZznaE0Vw5e+ehJl
3wY4+KqEZ3SZ8PAvDo9N4G1nx0E5VVYWH9bys50O53fgg6i1OKHWK6GcQZxKUXBU3B9aoYDsCZoG
59xph0k4+oydx24G4FgqAxxgTOJ4yZU+nzngRN4EwNnJ2+8uam71Iop6k0YaSMPbQkjDemPYKLo+
6mwW7LlsKwc4gey0Wlhf2FLOGk3ep/6hze+Ne+zPpP5YOj5W8VcraTH/GNG5H63fbjS6RkhY9GpE
qXW20AWkr7HdoHbAYJkbHYuVBO4cJ2l6wUDXOL+sCfwc198Rr55thN3mxWqgDwUYk0ZBb9LbGlCF
iW6cflzfO071WXileMOAHh3845O54vt0XEVSB5LbMSpFCk6216g+WozQXJtSUn3F6qotR7QZ3enD
eJrc3G0x6H7zD54qcpuJHqvD5YzDghCTlG754uY0gjPWrEx8XrXpWbEZcBvlV3kq8Yb8aLg0I1Tu
L1FAO6Y6DvmSpwCVtuTp9xFo1NI32JTBO/FZC3iro7Vg+UZ3BbDvAAddTMSZ+higzBjbJ3zCMSm1
Xh2PsMGkLvYqocEJKbdw6yKyxO3sZB7KEyrOf4Rv1JxMJhZvDkMJUpL5EgioSgiNpkHXNtZ750xL
xYHv1valwCVBwoHF6SPx9SNya3YN1c2IIa+maz71evIV1EQybBZupDrdlIx1UZGKxmrLVbYmuELy
DAYCxlj2n7mgPJo3UY+C/2EWcJH8eU2lLoP9/OSw16GrSlkrPWC5j9i5HRVysrdUMx18kXfKupCv
rnRAMQ63EvS2acmYh9msXRpWQhWidjetDVP6TndXQ7LeDejp9HSMIOo8AAAgE+OjOCgSgHssVHNk
fFvnSWhyZSVyckLG2LxOxoPLHGGDqGcHDfRohhUZAa3FLwsLugxKyoqzoi/60PKp7st6YWJAFbjO
IK5hurHPyJZ9FLsdYvHTLLBgRHNXBj3o30dtMl6rS/v64okaz3DJc1ZlA6Hn/4YOw7WVGbzTaNNt
IlNet1SmdpriYaJ+L1ysM2CPRkbpKyoSVnDri9wl7KJE8nuLbb7A5jpmTjv1QNWt15LUk+ztfQfw
Ulyq3bw+GQxD7gpjWE5j13pbpQ57XKD86hNUSnj7wPL4JCGxfbFDrDD3mpuFPkKTZna+Z9bMmzea
1fgIwzE214BjUPQ0RxDgYi1ebLbgwF26hrfGsYK+YF251Wfh6nw+a5hdtm8YxrHOOSczVJtDn+Uk
8zK2e+h16lZ1AoIGVFUkS/6svOxqLGS6vErYR4YgoRHGggMtrvrjAfkcaBt37DqP83OKm96BLeui
7iDL7EHWLfVR0F+bEOcUPudNG+86deN7punE35ZeJ5KtjbJcgNhsCFEySzHcC1fjaABD7YbBkt1p
X3+CkyrZkj8MKchOIJbpAFSMmfit7ZcD0+RMe7NQlZTK1nSz1ugJ3ALmSRPm/5H8oLueRB4XHJV2
Za8syayqwJFNR4mCqMk9xzb6swmTSDqmPWYXTfpYlcy6JDE4cMu/Wsr2LDe8ESx1AOoumCJGYzbq
eYfgT+dwrX1N+mPG8R7EwwvvQe3XksmKg1cpiOsPw8jpkCE/lxHtwOr4xai/A2J1Qhg8wlFhh/tF
ayYk/NpHE93eVZGRkfSrSxkosnX7sP6PXlBf5J3c1Bx556S4F2XciTr1bATgv73u2z48B/CL6X+D
+LdshS/9fmNw3MiwZ73bxnisOlfFnWI8WR3f5u4kghLXgMOrpj9vsv+YyggPV8nrMS19Dl8bG7PP
izA6+N+1NiLmjP2DDyDLNKIZjDee8JwRVOw4r9tl6hR8bGBwDZxD8QYTw2+AZXrzSqSsdIEsIqba
sHWAw1MweFHAqPsBkb2d1AHD25mnSXdEoqSVID3dQRsqFz8t1XiZJQ4x6mHhu2FuO9jxmKKOHhAq
xG2vQ5AMRNwabZv3BeGT7Qb4SkPT0UuAvxFGLzZShnyYEfvG3qHSrWx3Qi5+mVLOTnYMNNr5y/pa
zBeTtVIao4ypvGDgeLQr262UKXDjzfZYbteCSP2SPCtN0e7WNdegzdofxJuHQK8VGWgyn5+QseqY
G6PD31lDzxIN0TV1DQsQU5rs7yWayRulVgGIDzqJguFgNe0XBqenTG+7Xl88CTETjyZCYGqSJh65
QFnZ8VBpFikr81A5QIMNIsnCz/VGG/qQ2qmGP0gnoNnjhmT6M2VyXDeymlzuH8UejArpOfd6i7nY
jm3TmlDOudu/2QZOgxSV/a+7LSjz+23QTN1yGhPIFakJkV9DryDOPAwP1clfyWbH4WdkNzE4p6L0
66M3DMT8ErIPI/63yJ0J/wwXYyL1aaFzYpunHWYXXgeRCQlScQzfhLSzoK+Osa2CgvmrV7XpkEP0
BSJaXzIOBU8BCYry3VfnJIzXfuWa3UBq/BkOfnYXKoh3Uh6j4ltr7+EzmDwbJjMDuhc0UNasvPAc
d19GLOhvLewCaGplX9rJ5kChLXpccSs0WnKwh3Og+zt98fM6fYY2zN0GZEVUOUwA08G1mwSsBrwH
v3DmsdCrsFKBl4wRZf9NQYMv4tcDFUfTtsS6YNOC8Imz05OvF6EplKifKdArRKJtrTTVCn09m8Mk
IYaTsa+VQXOY1SV1ge6eAFvOC7a3x6UuZ3kIRnEFWF7wDKLeXv3sVkOaSilVL8AcUgd9dGu76Fz1
cnrJFNnuI3X6RXkrHrRiomvxd8+hOuQ20esepbrVPHcaAwQGzceWqrkzOsZ4/Uu5DwFEmgxSxUW9
JnBGaSu8FkCtvlrTDmoYRP3VNLyg65RQ5fpMsmy9mpKyNrTP3Bqoj7IpP02XZ09+oqzeY3KnqmX0
JeQG4pktwZt1NChBond9GQX1a8mKU8wHJ2qzjN77TMMbFW6vC56CUoppSckS3KeVKVRjUcMfwHGT
ARKt8RVPYy5g64e5kBL/Z1aJ9GR7CJtpCDNCZPcf4Ctkhn7uiM1owtOG3pi0Xt/LOgCr6ptV9jpg
Nsnh+gIuO3D7taLhgOMU4bjkQ6WfFKwf0ArJ7qTlx+4wcJXwYsGekMkxT4m7hE+glIoLsOFttTIp
bGzwIIPJ06Nb/4ZBX327UPrHg8/oZuRNo1zgYVFfktiBThkrBb+8kj+OBBK0Eqq2Uy1GJwtGGCl6
4LHxd83NH5PofAsy+14xs8vlZxudiMv/PCwYUFQBTGLJ0FX8wBnBBXIE8CKFffHJhHdKgT9+jmx3
w0ctUjScrquW576A4fvR4DI8LQ4mwqNqvQ8/uod++LklD1+gJxpk9gJVVHZg+NmVRYPMa4YBe64X
VpnT93xs6gCmikKhr/s4JIDJzukYpUK+E58wbTuyD3C2l0YagC3uZunDbcPxh1lufyEJ7OqNkKxx
TBU2BkXdufZ/ucKiTBFc4vy6aaiY5bB7O+LlS0Ns4PSWknnwS58Pf2eDMDVCdFgz48h2nSXSC37P
u6GU5Xp0I5XhnoKedmK88Fq6gpcnjNp9Cpgzo3VVBPwxArv+0t+qGEQTEsVSk8cnl1Z5VGEEDfeF
WuQ1cjKrJZjyU1+JPKZ2wMbCY/LAupzo3nNOYxCFCS1bTvcOyS0PVlx3RSRZab9vKmuS2Pjzi4H6
vticwbIBTBLD3j+jqoPf9iqY1OrR39lUGT7HZ1M3gTpppLPWY3bUTqGDXcEOHrHuLDbwF2ywKqVL
CIwLC9ZU3ZY3OPD8fPF1h9ywgrtIwRo+q/beihc3ZOSz2uBn6n+ztQ3iVTXnTfEH60nmjSvjtwO2
DZwPXqKfdr50AeUGFqxDp4jieKqlt6R2wQQWtDg03w9enIO0R2jLMayFY0jCx7VrHBPiAycppgl5
N7wiPnNzuk7zXRIQoju93NNnEP9j3NTKZKv2VTOaarQ+jFYT0LS3hvpO4/TJmp4caKZcNFikcf3k
/vUNelmJ7lRZ4fPadcjOAn8ZoGlXQFVAeSNiG0vTidjaBZ9tFoJmZP2hBUbjyV+gfHRV9nYJPurA
wH3c9reY27wH9P7Rtugll4dDV9fqXz72meoNHVvjwYEbaQVTZJyhUrphwdqxxKB5Rru3mNyOVczJ
bkYZ1bSYKhKhVfVf1EdPa8EkJmYdu2IvimlHWJnoWWbKPfJfGyTTBlJ5D/hT624SFlhlHnsJSh39
toQPAb2XMYswkI1u0krzW2tirex06AxTy1SEo3RxQCusHe4no/pWXzJyGGMFwa4qkBmVTf3aiora
8Sd6YF9iz7fhRACUb8pCRDj4qLoSpT2iotf3u5oek8rRdlB9RkIFX6I+ja+SokzDWNQPQ15nixBf
0myb4ljqGIKAB05CcjHpk1wCjU6Atk1nR5i01OFXqurmaFvvvkczlcgs1HOA3Gm9tIOwEddFC5EV
TsNu5fF6VpD0oAjMiumkvLa2HL6XDqVkI55cHKOryPdQMA7x5qc4/Zcz+QhHz6Hu9+G4yPNa1khW
FN8//vRkwBU4xvclC1eSmkqYkApB82bJICP8dEGfYZw2Yl7T22aF0LSlG3dKLpBbRtJjRnfnR+dd
7AjscuF9wnmP5kbKV00fnkDGK05EJVVknzr5qwTMHUSyAugSCxy+rAbXav7XsqwCBjqaRVjM48Ac
u2SMlvwCawI+GT5L1MaAWLHDTgGHLFfcEQodoFYZN+myw/XXK71a2FdABnK23lOXgsNpmNPgy7WX
CyC01rCmJG5DNEvY6ECFi1Mpg81n/U8p8zFV6IqkOGkFKpWkLubrq8kUSSTaCitUMoOSuCf4DV6D
WtZkobQ5dafjH8TMog50yo8OH1mtczD9DsNWm5gcl9LCfpEK38cdvknjMFfk92+1sGooSjtamhOy
B1fpZNTk5dC8cokGhyflQDCr9hOHHoprYOa5NNF5iY/IMKlOvFcxoOaVpJiLyJfTfnYQuErqakTg
eArpTmiMK70WF0t2frQP8NCCbkfNNFkVHpPJ2GsOzFM1DsHXWbDIlHRglNOPzvU0Eu2qTzxBGoyA
UiMLmi0HwGyu/zAlnzBNImD6q6N95NymRI6u2pjplEv7DcVzTDK6ZRLlI45/ByR0WdRY35khy2UN
2HDrO7aKJVcOtgDkWWufKrebyGbEfLQyBmoapNnO9Sl1tusz03u28CVEZ3qAu19omKX7Dc6ywxPL
0O5kJYwiGjUdgCJXNK3rAJfJWnOWyKScJy75n4jTwx6IJMeKSlcYgDBGYkqDXFkAzKC93jAkW4XX
BRgfhTE17/cB6nyzOuWjOCft1UcihzgQAgJVf3Ikp6Q0yJu0qznnA91OODRnjbC/Y79gPs/N8TyC
EmwRQvnxPICeFKAbJdDQPjXsvtsj/6ggvBWHCvae+EK9Xo36tsABmXYCZJLc0pt90vGh3zZ+nJRI
Cg6OxMb3Ym0UTmjfh3r4RoFe30EkarBiM2ERoO0UwzO94/qdlJbAk5oD8dT5czVuG4h4MOIP3Ea/
kmp6PoljxJYeQVyTPnVreH1sT+OFOZ7zK+d5FZbRiq/9cGotnAYzBq/pv6FfivmSsnFEvADfrTYv
qNsvlDW0u5/Xwz2XYbrQlh+exZvoJ10I+p/c8UQrMWi+05YIpAzlQzfYw2sjM1B7REm4Sdwrqk/d
zdycvrSHW4BZp2lec9yfiea4cUbGI7kx31qGlm16MDca+BUtgZVzGQx5KDKHTsGZo4ynwgwee6X0
4v+XScHolfHz655UCAJ3IUjR3ZhXikn1O89ctOHkgBiBSBDTRx/lHf9dtYon58deZRV0IcypB80A
9laA6x33CZiOMvDGtcZKfBjKMGHtipYajScs2Xauf7ec/zFm33bg0ICRTTBN8Kb3E5/QNZeya4fI
erefOvAoz7J5pYlcq7RNe6gkmPBj/FMEs1oS9cQbUuMinleslS++a7MjesCzpp5TfWu3aVRcI54V
l1bDE+CXoKxXEloEw5eW0fGOuqykvOXuXoZ9NwYq8QqLfbfjOAOC9PJaRoXj59htlfvE2WD1nWAo
JMO8YEDRy42TTd36xStBNy4QihkDaJXMqUbEC+gd88qBSziNmAVQXeoyjjIyei5ZNYyj4zF7oYnt
JYlBRZdpkUC/SnEvKKLPq2sv/zmnhlnTPbfBkobdpM9Z66UzXKUWb+ct3abyJsuFdSWu3Sh2NEb/
AlOqF/TRxLO4BrsCvted5C/gSc/Gd5L0djdNS3MFdKbwfWIf01VFf+leY2Gq3FALSSg5LcFjb9Xm
hy8owYQAtZAqbPJr64O6uvOeNUj+orBkwXRox7NpFz61o3ogM+bDunye25Rg2YOkozMkI5gKYPI8
oJDOTpQN1EK4SY8ac4wqIFVcrPZeEz5xNgkrV4QKZ5FngFLEPRJfHgAJU3GCAXMueQGH5m+cFhiv
pAAT2WP+FkzgRAY/Wpgwqj0hqoaB9CW9VqTo5vG22WpCl1zUfbBqniEoaB2g4Hp4PvtLkjpjcpeC
P+3AtQnPEsPTkpbGdZfac+6iBl1CA6pgwJ7OT/HVUU6vD6gXMvwJQmtaT/gv4JCrKC3CMrmjHsrl
YQmFyUCXhZZQz4k9Vf1dxHKGb0//fL2NYucGI+WL40E6+KgArH3wHmrj1LCDmQx9HMYrkfJICuZv
5ezI0gXU8bW/OS6+DrrpslgnzyTk4JbVK9eqdZ+ne/6tDqPSZVw7dhBLVLrZTdPWqTeFtOWBmLZO
IoME6rIcHmbNbHAmpDvNsOif/UX/k+X4v8WExbwQSzz2s0hvT/QGd3d/U2eHuxe33hLsAZNHeEX6
T7CAGEvHij1ohFKlsQk80TsTZVr9LStUfRwewEPpY92W0EpQ15m1e2z6DcYP745M49+ynHfm+5no
Zy3jG8WvOmDXPr/EEN0NnBUp+u3U88CIV6tWEd76OD9ICT5YcDCVOo0rZmhecaWHbFWfJrmCTdTI
olPexBBUzNWTgLmoeHVDwMGjOwyMJAPcPuEqHdJVNoZSF64BWKAdne3d5Z3AWtdUYZDqL2Glztn6
UTTW2QgEa9K9VhMBVCQrKUltb9sJE89ZjUtpR+GAjmBR0cHfks7FVcRQE0/OXbD9QwuzzPYAl61C
mB+WrtWnzh5eVgNjhBIOno2qiyFVeV0NerFoBivRm2xdwZ3hJgD1Egjr/Hx6I3CLcKm8kOXycBzA
CJVc0SNlivZ+yzhvT4szVax2XXjpP/Kh+yNZ5IuneJC4RrH0Fb0mqOgl/2KY1n3PEL0pCZPMRj2x
rG3Y1cgVV4FswJ9QKmOGHVZszeVL7pSlgLegMnLNHisdow0PdjoychsiI/jwOv3aBLfs1MJ3ywar
RdDqvWysqy2b943W0NSW0gBwhxovqE3R+GqnV1e8Om2MVJGkmvwWzPX4MZdUNxcmtMgGD6x0j0Dq
YGgZztNJEtckAmnxQop/kFUGtBDSSq2TeUGurBZ91lQR/uSGciyNqWUSKl/F8k0wewMv4CpenPR6
ySeqBx4jS1AGJ7Vk1S8/GbmU7+ADsen34KRwRKWS0FoDiyvExTNCxDceR+Hx43Z71CgYw/nRjzi+
y3CFbNKHRNi16t00bzH65l5drigoMGGGOlO0dr7eoSByuy3IDeBVaztbTrn8qbWODBcN82fQalPl
HF5pNR4CpBchk/BmVqIxNyo9zv2zkIhugyvkIly4vEDHJUB8wR6AO7MvyN1y+6jzxFS6eSjKxMu/
FN5k1Z/AGchiCDwVQDJcr5hjaN1h2W7D/88KrK8sPsVuL/sE++2maYHODFVn3rVT06+tnW1pW3Zd
e4ZyGj9b/uYQG21pYuPoXB92Np86y4CyEP8AeWpHSSQU21fIIaIOPRmB/oNp3XyuANfgEx/s1mTh
by/drrs85Foduruii81EQCZijVZbNMpkP9099miubJZAnSw6sOsiw5aBWCuOPNUC+hJXdQY4ochk
kGVaOLa5k1FMKEUA2VVC/yU4VS/cR3L+mxYIOFYwzWfaPhGxq04mriGTH6BP3VTxBsm8RYYKRIzo
dTgBiAPn3lFROu7ky5jURTnNq9a9wRVYvIG8MmbuRqchAhZMHO43ESWjHbdddJz4g6LlLlWM49Z6
1yCquZC9Sul5QPTIsFnZLvd8TLjje4EtzYi/GyZUrh2W5Ll/UXd4dSmhEuqVvRxvNg+vT7e4CGvQ
B9uiGiMMLNsGWUKYwaYqPpsGoheUSOWmMOSTn/UVKwDcVJpSWdJPXqTeqxY9PHIep3goTVdCj7T2
magjEudyIFzMBfHCGhzWg9XLj7dWkFoqPvfRb01k/m7ysMyFdyqoE8oykheXujCeuDI1nkB2ra/4
9EWPX/oXvnITmpkVuwt028mAOrbcAD6D0IdZo/msLysOECyvkefBpV9iodwi8lk8O8QqiCODwV6B
hJ4en9fAIeJOOqpgq6Mem/7jQ+d9CFXSCWzXsjIZ1Sg7eADh3SihFPhszUKV2HAv6/Vgy0nMqBC3
Og/ETVcFBu4CGpUSShBR2zicpsskc2I=
`protect end_protected
