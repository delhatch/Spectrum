��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J%�c2M���xWF�焲�b͠��ȾY��4�M�0���+��l��z'Đ�OH�2��K�O; �=��i������Z�H�6�P�4�\=}�XW� �cE{ądu�Qo5���Յ�b���*"z_�P�l��ЗTRE�ٝ{;x�誋k�'�W�~i�e9���˛j��&/�}��琕񺾾���d���<C�$�b%�qe����H&���R͹������<���l�p�d=�,�'P+��!�?3dI�����7텼8��4����rT���(�9C� g�p��`+Gp��}�%*�:q��m�j�u?��	�TJ��ܑ��=��yqh8c\ΊV}�Ss���;���Q��*��B�5U�׬���tJ@�;1T��-k\n�vr�'���F�`�ݨ�ƚ2��z�$$0�N�uʆ*�(�K���#uX{�%YY�zܱ���$���P�dt-L�w�kڎ� X�u�ZCP�	���V�G �&KAqV����EO��'� �r��3g�C�a3��)�q0}[:@�B�����7����zF���Ȋq�ᚒVˇ�q����ţd.��i"Wn��!�es앗6�y�����c��ռwꆙ��RD�8.��s���`����J�AvzX-��ǳl�����$�!�I�Ͻwh2�~#���%kA�P�F���M�+�yJѡ�7/l��gz����B�'��R������D{�#)Z{�R=��,�	>�f�ɔb��Ay�(.m���(����H�>C�lV6����^�Ք�H�|���U��T�F�WU���X��I���q�H!��1U1���5����+��,e��)�s��<V��{��{�)�]	HF�9HW��a`���mg)������Ֆs���D����=�]�	S���9��{�����v��Y���u�w��!`ޛ{�ڨ�$�z�_;�N%V��IiCԺ�Gv���
��>�i��� 8��E=�q}:�!tj(���e-��b-ÿ(3�+�\Gh������b�Z��eŭ�hx�(8Y�<V&�Ѿ��c�E�*����RY$6�ZV��-~Z�}A4P69���M~�X��x6���M�{\�E�hug-E^&��9�ذx��C.<���U ��iq��!Ym2O^
<R����Iր婢�G�iU�@��l���2([Rʡ���C�²X�>
j���Q�N�_N��V�=Q�>�P\�n���g�X�u���((��n�",�4�����q���Lt��;��~�k@�����$~8�Z��I��]���jRZ�CFA���l�|z�(V˧���c���BT�7�����}�f��6"O7�.������e�Bnq�e�!�H۬�޵lX���#m��.��&�n�D�$ri�L�����{�çC�����y�'p�����J߭`0~P�X;�1`oĳ�a�K?iL�]�!5A��³��������w!������<�w<Ѣ�^��X^֘�p�P��wG��0;��� z���IM���SN��Q�$�.�,k��\;t xHY����]1�˪8ׁ&ʫ��@���ʙ����ů��E�P��P3���z
���8�Փo2,�:��0@�1at�Qn��<��`[H��74��!}>TH��\f!�69*���J�ŨP=���ȗ�=���
}S��:���*|�`�8�r�5n�!�V��~�9�y�v�u0����vY�[�苭�D`h�FG��L�\6�K�l�8oX���%�����ZT����J�^*�׵R~〰G�����ޝyk�r"��饢�;ȆHaE��mEM"�A�|�t�A�Cλ�<����ؽd�)s�����V�&:t��e��cc�>a�c%�;���*�D��	�,NT�(���м�'P���;����|��ߢ#�*��'HJaak���m�����x�d+����n�V���'�|`�Q��S-rY0��T]�l�\�z�+�!�C̬e����X+���|�v�}����7\�-�dp߾Ӳ��K?��|�QCʵ���Q3��%��FӾ腈CD_c��:�v	w��"����&�p޽;����	��tC+���DH�-���u,0+n�b�q���ҧ���VJws�#�f\��&�I���F;��?�M-�d�.1W�3{d�aͱkeҌ�V�Ybk[2��>��r@R�&��.��j�l_�����P���0=��%����.�K,I�8.E���q��>���J<v�B�C�x��B�7�/���%��R�:,J,U���<?���͓R�g-�Tu=j[�pY��\�����v��*<hG��HC�pdi�|�����S���J�ŝ�>�F�n��'��`/�Ґ'`V�I`���"LX��O�Q���j%q>�������_����=J>��z�G`�aiEj�ˎ�i�A�g��Y����tu��o-��MQ�ʧ��b�1�-�C7�?�Bj4�M��'��j�[mK�pLa�D�vj�ϒ5B��@��ö��Td�?�`u(S������+�jP�� ��$ˇ��'�+*��HL��S�6��k�Ϯ�,-�h#(�옻�R0ľ}����+%�h�=]�j	&�������/݉�f���K��>��u��Ex{=u��sR�AuFsD�:B&D,u����G�N��OLDN��bk��E�}]�p�n^��DJN>ncb�)�C�W�̡Q�u�-^�n��I
��jkmһ�8�*Y�q�~�nw��p�]�C�"^��ڌg�:>0И�{��qҨ�܍�O�je�����)����ܺD0>.Z�ii������T��E�{��*cJ�?���G�7^]$�)�S�J��l��w�p��kJ�G���r1���7&N�m.����Fz���g�V�׮S�X���{�Km��F�7=N�15D]{���7;�0p��;HD�2�����K���ː����W�>�+�'��u�g>|���|ED<��'Z�5T820�؎]<2�B�L�8�
K���G����n��rVÙ���͌���y���r�5(����I
�\��!���0C�|��<��V���޹��7��ނ,)���	\s<�@'��$|�#�ަ*�]߼���4�%I������#������/�x���P��S�e�v��j��t����۞��G���}<L{12��)����+�+�)��TpQ3G]n�����¥�K7�mj�Uk������w_�$=A��^���=�-�o���|�v2�KI��P��]m�p_�z!�1��@��J\1����]�fń��Hc�� �|rB���c}�ѣ]M�j����"�}��p㋱�B����*9ru���s�s�QDY�� i����"��g�����o��h)ݓ_v!�k}C6C� 1�sD8'�s���0��cCD#�ofa�#X3��ib����J	�QY8��Ӯ@��j˓{��K,��*�����oXQ��k��&��{(��r�������+N���_��[�y/�N�$�A�b͙l4W�S�}5?b�ٸ�!�x�H���$`g�_��g#/E]0{f�<��NC�Y�,�I�E�>���)5�d'�C�Q�:�JeK5/́��vZ�������bAZ��4�-���7���¹�c�_K$lEU�G�g6��_�$�XTpDo��^�OC��W��y,QWi��J��l��<�M�v��{�������ܜ0~����CPn�.�4����7q�J�(�J|1<b0}��%�o4r
a��Ve�AT���v�>��s�����w8WX�"��M��V~�	by@Z]3k`π�ݼ'-��rq��`^�K�z���y�+I�Mv-$��">W[�{Y\�lҊ�mS�����I�ys&�"�C�3݀.!�	>�f*���A���[=@����j j:V-�2�i�Q0k�V�S&��J[��Z�7���74D��s��MX{�ɪ8
����+X�=�d�h~g�i��Qy���s����W�V��M��'H �7`�4:�r��v/~��As���ru!�/C�5d3�˦s�/Y��s5�)?]/����щ�O�D��($M�^4`�LPa0�]>����e��A$��.��IUi�)S�gI?��3�ё����a�0u���7�����y2Z����?� ܈� ����=������e}v��J��&Z�Y�*?$�XjB��7XS�&�@ԝSM���_����yW��L!J�����Iu׀�!���7��U2tք�4N�����2c��orkO��1��,5����W�f��{���E#[>��@E�����K-g���I7�nݙuh�Gƫ���� 9'~/wp������ǏkA�
�m�G�����+����4��N��5(٭�O�ك�~�M���Ӏ6�%���F�����i�}��M'ˇ�Nm�ʕ�|��04�fS�[��P��tR��AN�A�H/��"_��TI*�\d7$"��+����W���l�׮J���T?}|U��H)��(5��#�*�D;���,�8���S�*٧R\�޺IgΓy&&��K��6��)A}��4\D
'��#������eq�Л�3�M5ZcT�b�ܾ�w�f{����b��Q4Ǳ��1:������1`�Q�i�.7�ҵ�ͨ<wٲ?\s8��D.���"��^�85�x��GQ\����d��6����8�F -u���:ׇ0����o|rwo2��C>Rr!�m�g�Jx1ҽ�"w��"B h9<4EI�6�SW���&�Oct�YJԎ.H�E��o��G3k�G4�Gl1vg/ Q�Z}�-Kk�ئ�17p}��p@vA�H:Z��@�Pk��H<��2E�a�x��2�jok������xgƮ�N�8��z�B+�eu?�*�n��L�s a�#���Z���Pl������ݜG��T{�PSo��Tt4�o7.���(�jS
��v{�q�N��F���ar6/��H7ԁ/4��'���`�\EW�~Dm����@)�e`)&)z����u�Oo-�|��j�ϔ�0F�ݨ0\�@E���h�[`��f��A�Ck���������U�I�(�F��崱*О)23����A�LG�
V�}4W��mK�(�U,d"�FͳD^�G�l�� ���""}�=�WN�|`^Dg�l��xbf��!��n{�[�P|F����Q��������֏�&&�?�h�58@�������J5wG<���ca3�ҡ��M�~x��k�Zб	Kzf��)%�����Y��D�9�8�m�|����F�H��G'�#۟LRP]�_dH��S�5'>�5�Y��_F���S�dN�%_'�͑&	�Li�Y�5S�&����aGc��OH=`�PΒ����G"���\o�p�x��O  B�z[�=��
7Wd
�j��?8{0�������U�u�s+/;O2M�$l�d�,^��ж��|��e |�P���Q�@ge.�hcU��?r�ำ=����� Q���W����v�M����9����P;ɮ��FEi�N���[�����b=Y.�R�C�蚙w�L����D����*�E8B��g����^��K^��7��̀����3	��#^�zH����VMuRQ�?��Qe���81ю#�l@����>_���\}����=�~����ل*���������k�9,���s1N� ݞ,R@wz!n�����WB�_��v�<��Q��X���Vt�f�+�9СkG��@�o��@x�� �;6��V���Pү�&�}�:����y��;�"㨨�>rͦ	e����r����(��L�@�ճXb�T�����0��B�+^w?'\�*@��p�<q��+%S����]mfBƈ���	�.�0FD�&%R���� |#��Up6���2�/�gr^q�W<������3��55@���8�-�l�����F=�9�	#7���?�g�J�;�~�6D>�S�}5��	#@oN�Ad�D!p"[�ҳ�e�u���V�zp���ܼ2e�Y��c�x�����15km�xtIs�H�M!��HU�G���wj.�l�S93{�w�j$���1��kֽ�۽S|P_�o����v_Tsk������֓�"�󫱮(YO��i�M������L]��SOŘ�^.�O�Eۼ����+�~���_���W�B�Y��M����s-S#[P�I�5�������i�s^��% �û[�ɨ�˴"�ۛD��VBx:Q}���\��9_�A�h+�?�I'��N�}G %��-�a8EY���n}��>���5-�O����_������:ܽ���'|
�'YP.tɊ`�*J$�Xa��b��ȁ}*~nu�W���P@J��ŕ��?�э!��{� +�Cl�%x�_I�>�<m�s�Zя�;l�o�$��DT$��0d��/��g�x��%����}���'����!F4N'T&o�y��##��P}���L��t��q�-qF�lk�5���D�GQ�c�߭���������)�7ԫC<g��_~���
��*��p5�m���z%/���>��l����mV,J��^�Q�e� ��3���F-j.���S#�-7bW��-(���'ş�-��KV�a����(��y)���u�>�3�S^f���<�N��r�������%�[�-�M̖�w�f[��yO�ş���v�Sц����ˏ��u��яcQK�'��	~��Q�Lm���Ǭ$��vhn�s���YE�6����ϩ�����A�q΍LK:�\ƨ�W�6N���1���r|�'k�F^�����@���iRz�������,�`�&D~����F/�
�`X���](��.	���v ��bAmS��"S�BA(B�hz�:y_g�ت��;�57�)�����<�v.���y�-^
�yi���Grm���`�=.wt�D�h��*��F��f3-�pI��o�F�cڳ�O
Ba�r�<}�7�e;ʞ��k��>G�d{�3 �u�nf#q��>�
Et��K��W����4^Cĩt�0,Χ?�#�<|Z��WJҢ�����#�����*�����0[�5a/ʀ�� Vt�s���䲆���ʞ�)=O�%o�bP~࿃\,���ܴq%����]��k��$5]_�p�2�ԚY����mvU�E�P�B<��e���b�T>���s���]� �oBS�q�4fTfj�.!�Ny���B�x��)~�s��g��H�Uu\���r�BqE	�1J���Z���gW�F1�ǟF�d�7����g�A�� i��L��zy���}���� �P�Uw ��*Ohߌ�dB��j��Ľ�+J!T)�k@<+?w26sy ���n�|º�G�mܼmp�uv�}�<Ϟ���dg�a۪P?K6M�P�S���l6�n�|��?hK��O���͑)�S���(N'c�b��&j'#\��(^�D���2��p�
1�g����P��ӗ�Z�`�X&q��V�!���*ģ��k��m��*a�b~�
͘�J����uA�o>/��ހ�;8 g'��5��-n�q.H������,�ٓ�N����)�i�ɟ���fC~�Cb�Q�A�A������x�Ѡ,:Z�4��t�2��s�b�b�n�g��4�D2\ǿ���
Q��5Fm��{���¿��?��*��pt�|��X�Y��V+��X��_&f��$Z 4��\��l�h���[�x��6;x �y0����PC�\�HwD8��!�gސ���N�Q�t���磱�9�й,	L���ҳs�пkͿ�Z� ��%��9-�r��=�)��|�t���<T�ɽ<<�R�t�_�����p?�A�m��/bR�&H�kPl�_4�`��N��jb��Í�����3��:�N��� .�}0�:���*8�rB<�0��m��n�l{
�A9�K�^>j>�5�����裣u���8/0tL'�#�{�f%�_o,|�k���ĸ4����gެKa�x���b������"�Q���$t�I��&�P�{�֑����U�4G�]~u����nϳ��l�t;��d~/��'iA��:?T���@R�f���t�l�M����S�]�K�Ђ33c��� 9wW��>xC;�9��~�!�����;30	K`C���?��}����?˘|���������o�!L}?p�{}�<�)�����w�P<��S ��x����;���9�_u��	b��k��������טv���D_��|ڠ�>�5���Ӥ���ᗯ%�(n������0o������k�����A;��~Z?uzr�:�(������|)�������ܱ�OûWfW"D����8�D��v=�^x��I��"ҲLy�������E�Z��.+��ГH.6����y�P]|��*R���^R}�2��~�9�j	lwB�T���}黀Gr�WǺ�I��R�%ܹ֕)��6)Z|�\I^l'�>
�_�� ����%$��(qB����)c@�C�!�6�����C^��%��N6l�O�L���׃n�3���*[�x��� DZi��WJ�G(�|ϩ�m�5�
OA/��ʫv����!*��%H	�3����#fZ	߉��}}�R�($��K�	��<&�|x�ϥI�|cY)U�@���H0.������"W�xM�l�G��(;u���s=�j�/=� �gM�ӟ��`!2� ͎�}ŔM(2�zӠMY��؇[������8*���Dጆ럌'�f⿣�W{��[��r�����	�d�>NI˃�K�4�f)�U-dic�hab|�lHs|�Bcs���嬼���J��g'�ܷ��g���@��~0���G=^�����6`�fV�Y~���Eէ�e���������Y��?��B�N��$ff��'��{J?��Rd�%D<�+�ܸƌ��v���y���1����lG��ƌ?ߌ=I�q�^������`.�/T���u7�m�(�km6�Xbg2��@&B$;ގ�e��{�Ċ2�)�����(�be(���pi|xm