��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k*(\&��Y���z��;����1~;ó�!E7+ Uߟ �v��M�a�v���]�P9�Hq��;��p3��W�Op8>��N՟�8��i�yM�O6
m���h�V����_q�
ɏRa�H�g}�63t���&�X�~�^cȮ>�!����;R㿆�UHd�D8���5���_%� wt��fD��z��E?]Ck+������?�]�O�q���L�;�`��͐��wg����E��q���@ýW_���B�V�7�y�YݯŋI�Cw��9a��L��ݍK9�#�a�\����W���k�K�ٖ �gk{p��¸b����2+��Zq}�@�n���y�R��@_��U��`���9��e�Z2�XY�W�P�`�C\sq�C?�q�9K,IB���*��h�%�8��觘A$<Ȫ��9� SϾɓ�ۓ?����0�
�`�P���t�� GV\�|9��0�!�فp��l��˭�|�%����(`��1� ����
�$��U�^�pc�Ǡ�ܞ^���i���)vH�L�8c�cj]������_S_��{;�}=�D�-0*�kn_\U�{}�2\؄H�J22����
��q \
��N����?�_��6��My��Q+�����|&1^?����ڠ�VG��`Q�2�l��e7��S�"���"�(��U��������+�x�S[@�|-("����}��;��9�-ëy�'1���|E#1�+*|��c_����㞘
����+�z\���Otrrd�s��L%���d������C;��,���܈��k�l�3��)���N��E1����`�z ���,��)�F�`P����z�X+�`���)ߡτ��>��?�~O���<I��T����7���b_��B.�L��1iy�R���V���綤6��N��3���R�@�<���b���v|���v�����x�$m�U�Z��עnr��T��� zْD�7�$�w�;��o$���ߎ�|\�GO�b�%��3��۩4p�!�]u����T��<0�ķ˚�ؓ�e��@�L"�F��
�D��n��Y�A'z�q�C�"�Z����|# ����X��.AN9���xA��oa�Q[�<Ow�o�no��#�w�\,���C�}L*i����SD�K�}B�x��Q�pF���[�'|jM�^E:��*��C�������zs��x�>��}G/��ɫ�6c�C#���h��8�skrX���H�����F.D;��Q�����."�2�2��VLfn���E�)X��I�R���~rv���'�y"���B)*'��2
=7����U�^\a��JI<��B˭�Å�m��W|X��Ӥ�RV��c�%���z26͓��]�{d���9�B!cZ2�;�0��*�����\�w�7�u��,�a���F�vs"��d��f�8��\�%�t�_��IB�V���d��S[z}4�	����nP��W�e�r2��s��&%��0��8v;ݏ�O��19���O�n�6{�v�X������E2�0I,��������PA8��5rˠp�Kxֈ�@;	~�LT� � ���3�[-a�Z�ߡ\�?P��"aW����yT��pc�6�$Es`����s������1&Xӌ�<B�u&�7���gW�;|+>c2o'�I,M	��_����Oq"7R#| 'Հ[\���;ܵ�G�z?H�t��X�k�4T��Gƭ˸A()����*�%��gl�w&�y��AS���qa��� ��A%��f�^!��ܬ��*����
�f_����cmŤL`�s���ڸ!^zb[Z_��H}&.��jY]��tHNg{�|�&��w������:K�*�ƙNL~zz]/_N�R ը��ʜ���.6�ci�����{������'ݗ~�/e��y�8��"R;`m��?F�W�}�^ɞ@��
o�;M�R�	�c��/�ͨ�5$��&����s�ѶM��u$�*�Q�89�;F����|��s��� �(,c0)��qھ��"i�,�����o��z-�W���q�d�s7G��Az��4���"�#�O�#�A0k�@��
q�r-,J���/��`�M��"�r`�u^�����f�(�V�V�	��	:��:������{�~-Q�ւ8L�<+��IM����?
8m�W/�]H�L��\�`O+�j�Uyi�ӄ朎���{ñ#�m?/�bk�8>ږ���"آՃj#��N��K�cO���n��֮9�� ��㍅~�Tu�������h�<�?�
�wt2Z}P�͉}�Y�/luq1��;\���R}0XP�e;Q���/��-5Л"���hm�v��,w�ScY�k�t�<�I�AhV憒�4�IA�3�d�1�vo)���^���Eu6ڏ�"
��s�+2��PY�&�MSZ�B9��t������}��y���ٶ��4�Υ�Y:!��S/�´�i� yf�ar��+�-�kyM�1��|L���e����KwkX��-Jŏ>��e2��	��4��Y��[2��s�!&��݉/����ha8���<ʩx�P��ĩPD%J�aa>>��j���Ԇ
eK�t�������&��u!��l���Oi]�R:@�$w��>.o62�dL,SWb2"ԶF>s���]�&H����L=Ä�`�]<������.�l�0��s5�N�{TP�����=��/�,CcC{�4��.`���k��~)*hd��
=x�_a�Kx����%�)�Q��>�|�>p�
��Í�Pu/[�F-c5Yl��~ۮ��Th��(�&�1$w)^q��TnB��G3���C��3���֊]� ��mʯm�������J`V�9�lL?Z@�i�d��=���)IF�kv5�"�A�L�X�K�:�Q�vnd�YB��e�74�	C'�>��(ͶH��Ζ�����Ѽ��}�@nC��a��M g�@h����,�V���j3�&��5i
���	�7��Sz��������.*R`kܑs)��c��! ,��Zcd�ʖ��37�r����N����3`b�jo��b"Z�T~_���']�B<�q&%�&
Ʒr�X"E��؉��ǃ���*~L��S�jA����}Z%�I�2�Z�\R��Fk�]����D�?���]��6u�K�覢3��_�0�7�ԪEM^E���������e,".���Mu �f�q)�u�����avJ���pQ�A�!1�pi�5X/a�9 D�:�Tc=���l=�Ra��W���Ʋ�����a�0]�j�F�*�ݛ�� ��|�qPw���P�M�s5���x�y}���
 a��Fk�>'���1p�%i���ǵ	�iƹ?5E<�� ���(o$-��v��C������z�
��O����̓�F�)�D T�c���+��Ϛ8_�Z��Љ\���\��BW�1'�@�w��w��1��n[ŮdNUX s�/Y@N�h�K;ti�.W O���Ns3���sS|H1O��;oCn���r3k�@H��,��X���4��_��
m��8O!��DB#U[�o�a'���3͊���m�W nn�fg�/\� Ԗݥ88�m}ڗ��	gs潕�}J˂.t���w&W��?���#�E݁�U�NZE�ݠ��(B@g5ƽU���".�����=8$�"�%��$����E���/����+����l%�!�8��[C+<�7�r���*��g)�!t+�B�Q�����W	cN͛��k2E���y�P�/�D�U{U�����[B��>(}�	
���_exx�j�q�����2�-(������;�~��oT
��Q�祁#�׿<��>8җ��?,�$�'O�IL|���a:Y���F�n�� ǚ>����sJ�m1D�}�,���ʗӏcd�=�&�ľ���=8Ç��XP���ym��3�!o��!x��  $�kO�Sg����b�Nů�6!ԃ.��x������W�#?�3���V��J�����ƌ���
������G��u����OeV�"���ћ����㲍�r>.���|���g�уoS���?[���-�i&:
��꿫�^��-CU���;:? ��D���[Ȁ�3�RO���W�Ǣ]ϵ�GJ�Y烀.A�?zX���J`m�Y�&�( �e�[��������IM*��}P����;3�;�1-w��̂bNWͶh���_1N�lIՄ(*;	<m�q:�w|�냆0�lvSo$ֵ�S���]�Q�����tκ��{C�I�Co��)GC	}��Gw�o=�)e'�����fF���1��<ʞ"C�G�;��'ܭ�=�d��Kn	�AN�*�L4���'��}��̨݊�$tv�A�F{I���P٣�z�n�w_<U9���0Y^-\�z_�|���Y�*h��.�b_�n�9A������[�y�eE������k�F�=���\�?1�<�>G`���k�����qy@I�/~��-��6
YK����t'�64�x���{W�;=������J�,�:��+�,D^:# �2e@t���/㧡���g�=�r�눶[[h+Y����������$k����q�%�2j�p1V �0����	�"̈�}B����Խk?�����U�	���u4�`�7���%�p�~h��`̦��a>z:ZTu�m����7��Rg"���Z Cڻ
��1K��4���)�L>җ^p���ejI�N��>N����@%�� �J/PwX��ÐGr9��b�I�f>Va��n�=���w�FVӷ���C�hD������7%	���U�p�t��G���1��n����D���ڮk	i0�/w�BJ���W$�'R�ؑ�H�� ���)E���اz�����ؘ&@PL�'n���T��6~���� ks�J�Xj*S�Q��u��l`�J��HW6���	L��p��b2��`s���4�����ݯ�����RR��<�K����K�d�2[E�jW<�Fw�ض󦓨¶��e�܈���8�\�<c䪜�w̧�ݽ�,�[�=w��)v�2��ES��	/^�[U�yjm#��I9�D��Uu�gi*�|5��c�}�k?���x�ϋ�wW�Ie-/��X�E�vg�%�*�I�a!�xR�PY7P�y��.?�@��1@�G��(-Lw۲+�FNz!���ke�h���൚��CIJ�=+�D{To��u֧[�f����B�T�|���;�Q���*���l�ї?�o�����ʶE��̋��������|o�U�
�7���2�����l����?8S����P�.싕/������H�at�!Q�b/�۰��J��;�߻�7(�R2g�*�	*w}��I�VlJ�~�=?��O�;f@�����C����c��9��=�D%��%���w�5O���oS�Q�ƓW��IԔ��f&�ぎ������SU���+�;�x�pwj9+wDj�n#�Fn�X��)��;�d��*bq'���9D6�Xs�u zr����X-��t[�
w�ZXo���yO�����}�ڏ�e�k�1��ۼ�Pb�W�}��3Lƅ�#���B0����,��[�'���.�/1���G�KH�26���=�8��7l{��{��z�|�$���&��L6%D��m�
e;9N<U�!}����^f�8ϩ4ܤ��_�%�P�QaҮ󋗽� j&��Y��91��e���b�i�u�
I�6c�7�i0�θ�b�R��`��>3V�#�ƏB�]ޥ��7�On��������%B��@?�I(Tؙػ�뷣�޺�QʬKѬ� $��.]O�90L�ܚ[�2�^��ڢ�h��V.	��v����Ʌf�W��f�A��H_	I�Q?Kc̰�]�0'��B�\M�fQ_$tԇG1�@�#x.����9'�W���$�gR�u���C��|����=����ڥ�7Xb�K��T0<,�d�J��(`d�;�&%���l���1��w֙�`9]�oq����E�ԝxR.o�˨���%��د�[A��M�}�RM-\� �wDg���#�P�IT�C�!���!�|��`��O���E>5`O^uj��;��1�l����,�!֓O�IR�K�O����c��~�|Q���~8��T<)�*��%�93��=	*����b:z>	ꡔ�X~�j�8��J4�}PӁ���Թ��O������Q�=�Fh37��8\���g�F��h��'z0z��a{3;Nh�jrT)7�,�t*�� ��� ����ɬ������w�e�8�1�3q2�Y��f��@eu{P)�r�сUQ�}{J>��{������܈�Gޖ��'�}��������NF�%����@^k�0�����s�8��<�:��_�"I�/#Y��$�
,珫�*��ڬbyG�\�D�W�7���D��C~ҥ~v9���'8&*��
^�}k2�O�ߝ8�UYoQ�,B AW)%G�b&�WxZ��ǀ�����8?��{���3����;��g�`�ϱ�Gz�m�ӹ�vc�����)�bc��ϩ��Wh)��Q7���A>�����A	�M iFK��&A��v�x�#"�6��5�q�-�m"a_�\�f9QN��d �J�.�(l���̼�C�C�\�[~�#��"4KL��G�����6.��LQ�Q�ʹ�[��/�zP�;��	�n9��'�r���y(G�������z��Z<�&��8�i�9�i}|<��������A�v���;: