��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�kT��!`��� Z9**ul�T`�;#1͆<A���W���9��߻��Sn��nh��]�{s!�7E�o/dW�'��C% �B�_�	�S�a�o-J�4|ȍ�r�hƾ�A�g��5	�F�āF#��se�	��QP�w 4oH�H���D	�O���J]�K���[�VU�a�gx0�Ta�^��H��.��ݝ|�c�s��M�g������.{��$��M-Γ6=�Sⓔ�V�nvK�r^&����J���=ɫ֚;�p������׈r/IK�h1q�5 +�b'_���v;��w��w���w�oS��]T%m� N_s��W�)�?\-D�6��{�_���&��Ԗm#N�7:��^ѱ{L�E4 *RߴV�7BL_
����v;6��F�T�JG赫n����iHna�<4a��{'"E�U ���{$e���tFܸX{�u�.��/�lr(�d�I��7^p�Aq9G�[���y]�Hi���<D���3"jM�⿵c�Sy��;&�����b�c����z8��F�j����z~��>���?h������J.7��J�**��t'cG6��)���@E���;�xd�7 *'U�I�U���\�:1����j'��c4<��4P2���B��I<:۬KRE�_��Q���`�ҟ��[#�/�G��uzd���.��w�����R|��?ʹLָBb!*�)RZr֚���9�x�����R?�,']�S� ��1��gLB��c��xC�YOʄ�L.)�;��H���G�شj����aL'��i��w��9@�ުk����WR���m���򾖣o1�F9m�P_I���_Ҁ{��d��j+��K�q�*��O�z�1+